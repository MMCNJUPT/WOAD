
module gemm1L (
    input         clk,
    input         rst,

    input  [7:0]  addr,
    output [47:0] data
);

reg [47:0] out;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        out <= 0;
    end
    else begin        
        case (addr)
            8'd0 : begin out <= 48'b101100111000100000110101000001111001110111100111; end
            8'd1 : begin out <= 48'b101101110111100010110110110100111011010110011111; end
            8'd2 : begin out <= 48'b101110000010110000111001100010011011000010100100; end
            8'd3 : begin out <= 48'b101100001010010100110000000001100011001000101011; end
            8'd4 : begin out <= 48'b001110001101111100101111111000111011100101100111; end
            8'd5 : begin out <= 48'b001101111011110000101100110110001011001011001011; end
            8'd6 : begin out <= 48'b101110001011001100110110010011100010011101001110; end
            8'd7 : begin out <= 48'b101100010000000000111000100100111011010010000110; end
            8'd8 : begin out <= 48'b101011010100110100110111111110101010111100100001; end
            8'd9 : begin out <= 48'b101110011010000100110110001111001011000010001101; end
            8'd10 : begin out <= 48'b101011111110110000110101001101111011100011010111; end
            8'd11 : begin out <= 48'b001010010100101010111000010101001011100110100110; end
            8'd12 : begin out <= 48'b001000010010110010110010001100001010110110110111; end
            8'd13 : begin out <= 48'b101100100001100010110001101100010011100011000001; end
            8'd14 : begin out <= 48'b101101001000010110110011011001110011100100011101; end
            8'd15 : begin out <= 48'b101101010100010010110001110000011011100101100101; end
            8'd16 : begin out <= 48'b101110000001001010111000110101110011011110001010; end
            8'd17 : begin out <= 48'b001110000001110110110010001000011011100001011000; end
            8'd18 : begin out <= 48'b101010110011001100110111110101111011011111000100; end
            8'd19 : begin out <= 48'b001100110011110010110100101000000011010000110110; end
            8'd20 : begin out <= 48'b101100101110111110110100111011000010100100101001; end
            8'd21 : begin out <= 48'b101101100010001010101111011110101011100101101101; end
            8'd22 : begin out <= 48'b001101000011100100101010101010001011100100001110; end
            8'd23 : begin out <= 48'b101101111010000010111001010011011011011010011000; end
            8'd24 : begin out <= 48'b101101100111001110110100001010011011100001110101; end
            8'd25 : begin out <= 48'b001110010111101010111000001110101011011000001001; end
            8'd26 : begin out <= 48'b001101011011100000101110101101001011000110000101; end
            8'd27 : begin out <= 48'b001101111000100100101010111100010010110010101101; end
            8'd28 : begin out <= 48'b101100010110100000110000000001001011001001111111; end
            8'd29 : begin out <= 48'b001100110110011100110100001110101010000001101011; end
            8'd30 : begin out <= 48'b101010101100110000111000011000100011100101010110; end
            8'd31 : begin out <= 48'b001110011001010110111000111000011010111000010011; end
            8'd32 : begin out <= 48'b101110001001111100110101010010001010111010001001; end
            8'd33 : begin out <= 48'b101101110100010110111000011101000011100101110100; end
            8'd34 : begin out <= 48'b101101110000011100110100110111111010111000111100; end
            8'd35 : begin out <= 48'b101100001111100010110010100010101010110011100000; end
            8'd36 : begin out <= 48'b001100000011110100110111111110000011000010110011; end
            8'd37 : begin out <= 48'b001011001100101100110101000100011011100010110100; end
            8'd38 : begin out <= 48'b101100000111001100110100100101111010101101010111; end
            8'd39 : begin out <= 48'b001101010111000100110100101011000010011100100111; end
            8'd40 : begin out <= 48'b100100011101101110110111000110000011011010100111; end
            8'd41 : begin out <= 48'b001101100101010100110111101001111011011010011000; end
            8'd42 : begin out <= 48'b101110001000010000101000001111000011001110011001; end
            8'd43 : begin out <= 48'b101100101010000000110011001111100011100011101011; end
            8'd44 : begin out <= 48'b101010100011101100110110011110001010110011110110; end
            8'd45 : begin out <= 48'b101001011100011110110001000011001010100001010111; end
            8'd46 : begin out <= 48'b101101100001001000110111110010001011100000100110; end
            8'd47 : begin out <= 48'b001101010111101100111000000011010011100100001000; end
            8'd48 : begin out <= 48'b101010011010011000110110110111001011010000011111; end
            8'd49 : begin out <= 48'b001001000101000010110001001101000011010000101110; end
            8'd50 : begin out <= 48'b001101011100001100110000010110010011001111000110; end
            8'd51 : begin out <= 48'b001101000011011110110000011100001011100011111001; end
            8'd52 : begin out <= 48'b001101101101101110110101010001001011010110101111; end
            8'd53 : begin out <= 48'b101110010100001110011101101011111011010000101101; end
            8'd54 : begin out <= 48'b101011101001011000101111101001010011011100111001; end
            8'd55 : begin out <= 48'b001101100010110100110101010010000011011100111111; end
            8'd56 : begin out <= 48'b001101100111110100110101010101101010100010101010; end
            8'd57 : begin out <= 48'b001100111001010010110011010011110011100011001000; end
            8'd58 : begin out <= 48'b001001100011110010110101100010010011100011010011; end
            8'd59 : begin out <= 48'b101011111010110000110011000100101011010100110010; end
            8'd60 : begin out <= 48'b101010010111111000100101011011110001101011000101; end
            8'd61 : begin out <= 48'b101010100110011100110010011101010011100011001000; end
            8'd62 : begin out <= 48'b001101101111101100111001100111010011100000101101; end
            8'd63 : begin out <= 48'b101101110000101000111001100110010011010011000110; end
            8'd64 : begin out <= 48'b101101000010101010101110110000110010001111110100; end
            8'd65 : begin out <= 48'b001101001010100110100101010101010011000011010111; end
            8'd66 : begin out <= 48'b001110000111001110111001010101000011011101100001; end
            8'd67 : begin out <= 48'b100101000000111100111000010101100011100011011100; end
            8'd68 : begin out <= 48'b001110000100011010111001100011110011011011101010; end
            8'd69 : begin out <= 48'b001101011011100000101100100100111011010011010001; end
            8'd70 : begin out <= 48'b001101001111100110110101101011111011011000010010; end
            8'd71 : begin out <= 48'b101110000011101010100000010010010011001010011010; end
            8'd72 : begin out <= 48'b001110000110101000110000101000110011100010100000; end
            8'd73 : begin out <= 48'b101101111101111100110001000010110011001000011010; end
            8'd74 : begin out <= 48'b001101011110110010111000100100000011100010010010; end
            8'd75 : begin out <= 48'b001100010110100000111001010100110010111001111011; end
            8'd76 : begin out <= 48'b101110001101111010110110110111010011011101110110; end
            8'd77 : begin out <= 48'b001110001110111010111000111000001011100101010000; end
            8'd78 : begin out <= 48'b101110010101000100110001100001110011011011010101; end
            8'd79 : begin out <= 48'b101100000101110100111001000110011010101111111001; end
            8'd80 : begin out <= 48'b001100111001001010111000001010101011010111011011; end
            8'd81 : begin out <= 48'b101110000011011110110100110110001010010010101111; end
            8'd82 : begin out <= 48'b001110001110000110110110111110100011011011010000; end
            8'd83 : begin out <= 48'b101100110110000000110111101110110011010100110000; end
            8'd84 : begin out <= 48'b101011100011100100101100001110000011100000111001; end
            8'd85 : begin out <= 48'b001101101100000100110011011010010011000011111101; end
            8'd86 : begin out <= 48'b001110000001010000111001010111110011001001000001; end
            8'd87 : begin out <= 48'b101001101010110000110110001001110011100100100010; end
            8'd88 : begin out <= 48'b101101001100101000110100101010001011100110100101; end
            8'd89 : begin out <= 48'b001100001100110010111000111010001011010101010100; end
            8'd90 : begin out <= 48'b101110010100010110110101110100000010001010100011; end
            8'd91 : begin out <= 48'b101100111001100000101110111101011011100110100000; end
            8'd92 : begin out <= 48'b101100010101011010101111000010000010111101010000; end
            8'd93 : begin out <= 48'b101010110011001010110111111001000011100100110111; end
            8'd94 : begin out <= 48'b001110000101101100110100011110100011010100110010; end
            8'd95 : begin out <= 48'b101110011000101010110110010001110011010111101111; end
            8'd96 : begin out <= 48'b001110001110100000110100001000010011010010101010; end
            8'd97 : begin out <= 48'b001110011000011100110101101100111011100000101101; end
            8'd98 : begin out <= 48'b001101011001011010110110010111110011011010001111; end
            8'd99 : begin out <= 48'b101110011000101100110010000110110011000111001011; end
            8'd100 : begin out <= 48'b101101010111111010110100101001111011010001011010; end
            8'd101 : begin out <= 48'b101011101110011010110010010110100010100101000101; end
            8'd102 : begin out <= 48'b001011001001111000111001011011100011100011001001; end
            8'd103 : begin out <= 48'b101100011110000010111001011100101011100011110110; end
            8'd104 : begin out <= 48'b101110010100111100111000110100100011011101101101; end
            8'd105 : begin out <= 48'b101110001110110110111000011101110011010000100101; end
            8'd106 : begin out <= 48'b001100110011000010110001001110001010111100011100; end
            8'd107 : begin out <= 48'b001100110111101100101011100110100011100100111110; end
            8'd108 : begin out <= 48'b001100010001111010110100100111010011000001001011; end
            8'd109 : begin out <= 48'b001110001101011010110110111001011011010011100111; end
            8'd110 : begin out <= 48'b101101000111111100110010100011101011000110110001; end
            8'd111 : begin out <= 48'b001110000101101010110000000111010011000110101100; end
            8'd112 : begin out <= 48'b001100101001010110101110011100011011100101100000; end
            8'd113 : begin out <= 48'b101011100011000100111000100010111011011110101001; end
            8'd114 : begin out <= 48'b101100011110101010111000001100000010110001001110; end
            8'd115 : begin out <= 48'b001110000111110100111000100111110011100100110010; end
            8'd116 : begin out <= 48'b001011011110101010110001000111101011001100100111; end
            8'd117 : begin out <= 48'b101101100111010000110100010111001010111011100100; end
            8'd118 : begin out <= 48'b001101111110111010110010011010101011001010001100; end
            8'd119 : begin out <= 48'b001101010001110110110111001100000010011100011001; end
            8'd120 : begin out <= 48'b101110011001111010110101010111111011001010110000; end
            8'd121 : begin out <= 48'b001110001111111010110001000110111011100101111111; end
            8'd122 : begin out <= 48'b001011001110100100111001101000001011010010001010; end
            8'd123 : begin out <= 48'b101011111000011010110101101010111010111111000001; end
            8'd124 : begin out <= 48'b001010111001110010111001000010000011100101100001; end
            8'd125 : begin out <= 48'b101001111010000110110100000010111011100010011100; end
            8'd126 : begin out <= 48'b001011101110001010111001100000101011100011000001; end
            8'd127 : begin out <= 48'b001110000001001000110011110000101011001000011010; end
            8'd128 : begin out <= 48'b101101101110110010110011011011110011010101001100; end
            8'd129 : begin out <= 48'b001110010011100010111000000101011011001110110111; end
            8'd130 : begin out <= 48'b101011101111001000110010000010000011100100101011; end
            8'd131 : begin out <= 48'b101110001100101010110100101101001011010111111000; end
            8'd132 : begin out <= 48'b101110000100110010110101110100010011100000001100; end
            8'd133 : begin out <= 48'b101011100010000110110111101001001011010010011011; end
            8'd134 : begin out <= 48'b001011010001100110111001011111110011001010010011; end
            8'd135 : begin out <= 48'b001100111100111110110100001110010011100001000000; end
            8'd136 : begin out <= 48'b101101001011000010111000111111101011100000100010; end
            8'd137 : begin out <= 48'b101101100101100010110110001111101011100110010100; end
            8'd138 : begin out <= 48'b001110000110000010110100111001110011011001111010; end
            8'd139 : begin out <= 48'b101110001111100010111000100100010011100000011010; end
            8'd140 : begin out <= 48'b101101001001011110100011001001111011100000011011; end
            8'd141 : begin out <= 48'b001110011000101000110100011110011011010111110011; end
            8'd142 : begin out <= 48'b001101110100100000111001000111100010100111000010; end
            8'd143 : begin out <= 48'b101101110010111000110010110111011010010010101100; end
            8'd144 : begin out <= 48'b001110001110110100101001110110111011011111001111; end
            8'd145 : begin out <= 48'b001100101100110110101101011000111011011101010010; end
            8'd146 : begin out <= 48'b001100101111000100110011111101110011011111010101; end
            8'd147 : begin out <= 48'b001101001000000110111000000000011011010010010101; end
            8'd148 : begin out <= 48'b001110010110010010110011111101000011010010100001; end
            8'd149 : begin out <= 48'b101101011001100000111001010001010011001111011101; end
            8'd150 : begin out <= 48'b001011011011100010101010000000100010111111011011; end
            8'd151 : begin out <= 48'b101010100001001010101000001110100011100000101111; end
            8'd152 : begin out <= 48'b001100001111001100101111001110011011001010110110; end
            8'd153 : begin out <= 48'b101110000010100000101000000111010011011101101101; end
            8'd154 : begin out <= 48'b001110010010001110110000101010011011100100111101; end
            8'd155 : begin out <= 48'b001110001101001010110110011000100011010001011111; end
            8'd156 : begin out <= 48'b101100110110101100101101011110111011100100101001; end
            8'd157 : begin out <= 48'b001101111011111110111000001001001010100000011010; end
            8'd158 : begin out <= 48'b001101001111111010101100001011010010010010101001; end
            8'd159 : begin out <= 48'b101110011010010000101011111111011011001100100010; end
            8'd160 : begin out <= 48'b001110010001001010111001000111111011010101010110; end
            8'd161 : begin out <= 48'b101100001100111110110110111010001011010110100100; end
            8'd162 : begin out <= 48'b001101100111001110110000010111110011100010100100; end
            8'd163 : begin out <= 48'b001100001110101110110110100101001011100110010110; end
            8'd164 : begin out <= 48'b001100100100100100110101100000100011010000100000; end
            8'd165 : begin out <= 48'b101110000000110110110110111000010011100001111001; end
            8'd166 : begin out <= 48'b101110001001101000100111111111100011100100011011; end
            8'd167 : begin out <= 48'b001110010110001110111001011011100011100000110000; end
            8'd168 : begin out <= 48'b101101111111000000110101111000100011010010100110; end
            8'd169 : begin out <= 48'b101110001010001010111000100000111011001101111101; end
            8'd170 : begin out <= 48'b001011111100111010110100110100110011010011100100; end
            8'd171 : begin out <= 48'b101100110011000100101000010110001011010100000110; end
            8'd172 : begin out <= 48'b001110000011001010110101110101001011000101110111; end
            8'd173 : begin out <= 48'b101110000100000110101011111100011011000011010001; end
            8'd174 : begin out <= 48'b001110010001000100110100110110110011100101001111; end
            8'd175 : begin out <= 48'b001110001001100000111000001110110011100000110010; end
            8'd176 : begin out <= 48'b101110001001000000111001001110010011011100001011; end
            8'd177 : begin out <= 48'b101110000001110010110110011100011011100000010100; end
            8'd178 : begin out <= 48'b101110010100100010111001010000111011100010011100; end
            8'd179 : begin out <= 48'b101010000101011010111001001010101011011101101100; end
            8'd180 : begin out <= 48'b001001110000010010101100010001011011100011011000; end
            8'd181 : begin out <= 48'b001100010101100110110010110000110011011111010010; end
            8'd182 : begin out <= 48'b001101000011100010110000000100110011100011101101; end
            8'd183 : begin out <= 48'b001101000011110100111000001011000011100001000111; end
            8'd184 : begin out <= 48'b001101001111010010111001100010101011100001111001; end
            8'd185 : begin out <= 48'b001101111011111100111001100111111011100010101111; end
            8'd186 : begin out <= 48'b001101101100111010110110110010101011011010011101; end
            8'd187 : begin out <= 48'b001101110110110000111000001100000011010110101000; end
            8'd188 : begin out <= 48'b001100000101001100101010100111001010111011000001; end
            8'd189 : begin out <= 48'b101010001101110000110000001001111011100101010101; end
            8'd190 : begin out <= 48'b101100001010011000111000110011011011010111111101; end
            8'd191 : begin out <= 48'b101110001100100000111000001000101011010000001100; end
            8'd192 : begin out <= 48'b001100010011001110110100100010111011010111111010; end
            8'd193 : begin out <= 48'b101101111011100010110111010001101011100011111011; end
            8'd194 : begin out <= 48'b101011100001101110110111110101001011011000001110; end
            8'd195 : begin out <= 48'b001010100001011100111001011010110010110000110100; end
            8'd196 : begin out <= 48'b001101010010010010111000100001000011001110111000; end
            8'd197 : begin out <= 48'b101100011011011100111000110101110011000010011010; end
            8'd198 : begin out <= 48'b001100100111101010101110011010001011011101001100; end
            8'd199 : begin out <= 48'b101101101001101110110111010111000010100010101101; end
            8'd200 : begin out <= 48'b001101000011110100101010100100100011100011110000; end
            8'd201 : begin out <= 48'b001110000111101010111001100001000011011100111000; end
            8'd202 : begin out <= 48'b001101100101110000111000000111011011010000100010; end
            8'd203 : begin out <= 48'b001110010100111010110101101011000011100011000110; end
            8'd204 : begin out <= 48'b001011110111001010110011011100111011010000100100; end
            8'd205 : begin out <= 48'b101100100101011100110010010110110011011100000011; end
            8'd206 : begin out <= 48'b101101010001010010111000111111110011100100100111; end
            8'd207 : begin out <= 48'b101100100001101010110100111110001010111100100011; end
            8'd208 : begin out <= 48'b001010010010110100100001100010000011011000111100; end
            8'd209 : begin out <= 48'b101110001110000010110100001011110011100010001110; end
            8'd210 : begin out <= 48'b001011010001001110110000010100100011010010011111; end
            8'd211 : begin out <= 48'b101110001100001110101111110111110011100011100110; end
            8'd212 : begin out <= 48'b001010110011111000111000010001111011001010000111; end
            8'd213 : begin out <= 48'b001101111100010100101101100110110011011001011010; end
            8'd214 : begin out <= 48'b001110000010000110110111011010001011001111010101; end
            8'd215 : begin out <= 48'b001100111010110010110011101011101011011101110010; end
            8'd216 : begin out <= 48'b001110010111100110110101110111101010111011100011; end
            8'd217 : begin out <= 48'b101101111100110000110100011101101011010111100111; end
            8'd218 : begin out <= 48'b101110010100000100110101011100010011100010010001; end
            8'd219 : begin out <= 48'b101101101000000000110110010110110011001000110110; end
            8'd220 : begin out <= 48'b001110010001011110110011100110000011011000011101; end
            8'd221 : begin out <= 48'b101100001101011010101101001000100011100010010110; end
            8'd222 : begin out <= 48'b101011011001100110110100110001011011010000011101; end
            8'd223 : begin out <= 48'b101110001010011110110011100001001011010010001010; end
            8'd224 : begin out <= 48'b001101010111101010110110101111000011100010000011; end
            8'd225 : begin out <= 48'b101101001100010110111001100001101011011101010101; end
            8'd226 : begin out <= 48'b001101111101011100110000101001100011100001001101; end
            8'd227 : begin out <= 48'b101110001000001010101000001101111011100101100101; end
            8'd228 : begin out <= 48'b001110001100100100111000001001000011001111110000; end
            8'd229 : begin out <= 48'b001110010110101100101110000110100011100011011111; end
            8'd230 : begin out <= 48'b001110000110000000110101111101011011011101111111; end
            8'd231 : begin out <= 48'b001110001001011110110011010010101011000110011111; end
            8'd232 : begin out <= 48'b001101100000100010101111000011111011011011001110; end
            8'd233 : begin out <= 48'b101100110010011100110101001111100011100000110011; end
            8'd234 : begin out <= 48'b101100110101101000110010010000001011011010110000; end
            8'd235 : begin out <= 48'b001110001001000100110101100010010011011111100110; end
            8'd236 : begin out <= 48'b001110010011001100111001101001001011100000111110; end
            8'd237 : begin out <= 48'b001011111010111000101101011110011011011111101011; end
            8'd238 : begin out <= 48'b101100100111011010110101000001011010011100101000; end
            8'd239 : begin out <= 48'b101101011110101100110000110001101011100110000101; end
            8'd240 : begin out <= 48'b101101101000010110110101100111011011010010111111; end
            8'd241 : begin out <= 48'b001110000111111110110100000011100010111010111000; end
            8'd242 : begin out <= 48'b001110000110111100110011101111111011100010111110; end
            8'd243 : begin out <= 48'b101011011101010100110111010011110011001001011100; end
            8'd244 : begin out <= 48'b001110000011000110110001111101100011010010010111; end
            8'd245 : begin out <= 48'b001001010001110010111001011101001011100011101011; end
            8'd246 : begin out <= 48'b001101000011111100110001000101010011011101010111; end
            8'd247 : begin out <= 48'b101011101010101000110011010001001010111000000000; end
            8'd248 : begin out <= 48'b101100000101110000111001100101000011100110011100; end
            8'd249 : begin out <= 48'b101100011101101000111001100101110011011011111101; end
            8'd250 : begin out <= 48'b101110010110000000110111110100011011011010000010; end
            8'd251 : begin out <= 48'b001101110110010010111000000000011011100001000111; end
            8'd252 : begin out <= 48'b101110011001010100110110110010000011001000111101; end
            8'd253 : begin out <= 48'b101110010010010100101000011101000011100011101010; end
            8'd254 : begin out <= 48'b101110001110011000110111001001001011011011001000; end
            8'd255 : begin out <= 48'b101110001000101010100100100101001001001110111101; end

        endcase
    end
end
assign data = out;

endmodule //gemm1L
