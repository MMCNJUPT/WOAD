module gemm3B (
    input         clk,
    input         rst,
    input  [6:0]  addr,
    output [63:0] data
);

reg [63:0] out;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        out <= 0;
    end
    else begin
        case (addr)
            7'd0 : begin out <= 64'b1010010001100011101001011010111110100010010010101010101101101100; end
            7'd1 : begin out <= 64'b1010101110110011101010010100110000011001001100110010010011111010; end
            7'd2 : begin out <= 64'b1010100100111101001001000010100000011100100110100010100100110010; end
            7'd3 : begin out <= 64'b1010101101101010000000010111001000011110001011100010011011011101; end
            7'd4 : begin out <= 64'b1010100000110000101001000010010110101001010001011010010001100001; end
            7'd5 : begin out <= 64'b1001110101101110100000001000000110011011100101110010001001111010; end
            7'd6 : begin out <= 64'b0010011011111011101010011000011010100111001001010001110110010110; end
            7'd7 : begin out <= 64'b0010010100001110000110000110111000101000000110101010001001111110; end
            7'd8 : begin out <= 64'b0001001011011010001001000101011110100010110110011010010001100011; end
            7'd9 : begin out <= 64'b1010100001100010101001111100011010011101110000100010000111000010; end
            7'd10 : begin out <= 64'b1010100010010111001001101110101110101000111001110010010001110111; end
            7'd11 : begin out <= 64'b0010010000101100101000010011110010100001011111110010100011110010; end
            7'd12 : begin out <= 64'b1010101010011110001001100001001010100100111100101010011101100101; end
            7'd13 : begin out <= 64'b1010011101011000001001010111000110101010010110111010001111111110; end
            7'd14 : begin out <= 64'b0010101110010101001010001001000010101010000101111010101000000001; end
            7'd15 : begin out <= 64'b0010011100010101100101011110001100101000110001001001100011111011; end
            7'd16 : begin out <= 64'b0010101011110101001000011111001000101000100101101010000110111100; end
            7'd17 : begin out <= 64'b0010100010101011001010000110111100101100011110100010101000011100; end
            7'd18 : begin out <= 64'b0001110100100010001001101101001110100110000100101010011001010010; end
            7'd19 : begin out <= 64'b0000101011101000001001110001111010101001111110101010100101001111; end
            7'd20 : begin out <= 64'b0010101101110110101001010101101000101011000011000010100111111111; end
            7'd21 : begin out <= 64'b0010011110011000101010110000000010101011001011001010011110010000; end
            7'd22 : begin out <= 64'b0010010010100100101001110101000010100100100011111010100101110001; end
            7'd23 : begin out <= 64'b0010101110110010101010010111111100100000111000100010010110110111; end
            7'd24 : begin out <= 64'b1010101010010111000110101010101100100000101100100010101011100101; end
            7'd25 : begin out <= 64'b0010010110111011000110101100110000101000010011011001011100010100; end
            7'd26 : begin out <= 64'b1010011010100010101010010110111100100111101001001010100001101001; end
            7'd27 : begin out <= 64'b1010100011101010101010000111101010011000101000001010010000101010; end
            7'd28 : begin out <= 64'b1010011001000001000110000110010000101000100000011010011010101010; end
            7'd29 : begin out <= 64'b1001001011100101101010001010100100100101001011111010101101010110; end
            7'd30 : begin out <= 64'b0010000101000100101000011110001100101011101000010001110100010111; end
            7'd31 : begin out <= 64'b1010100110111001101010000111100100011101001000101010100001000110; end
            7'd32 : begin out <= 64'b0010011100010000101010101100100100100101000100110010100110110110; end
            7'd33 : begin out <= 64'b0001101110111011001010011100000000100001101000001001000101010110; end
            7'd34 : begin out <= 64'b1010101000000011001010100110110100100011011000001010101010101011; end
            7'd35 : begin out <= 64'b0010101110101100000110101100100110101010010100100010101110100110; end
            7'd36 : begin out <= 64'b1010011110110010001001000101001100101001101110011010100001001111; end
            7'd37 : begin out <= 64'b1010101011100100001001110001011100011101000101000010101010100111; end
            7'd38 : begin out <= 64'b1001110011111011101010111001101100011110100101010001111110111101; end
            7'd39 : begin out <= 64'b1010010010101101001001110111001010100100010001001010000111100000; end
            7'd40 : begin out <= 64'b0010101010010101101010001010000110101001011110110010011011011011; end
            7'd41 : begin out <= 64'b0010101100101100101010001010000100101000000000111001100110110010; end
            7'd42 : begin out <= 64'b0010011010011111000111111100000010101011111011101010011011011001; end
            7'd43 : begin out <= 64'b1001110010101000001001000101000110100011000001000010100001001011; end
            7'd44 : begin out <= 64'b0010001111010000001001101010000100101001100011010001110000101011; end
            7'd45 : begin out <= 64'b1001111101101101001010110010001110101011000010000001111000011110; end
            7'd46 : begin out <= 64'b1010101100011010001010011110111010101011101011100010101100110111; end
            7'd47 : begin out <= 64'b0010100000001111001001100001111010101010000111101010100101101111; end
            7'd48 : begin out <= 64'b1010101110011011101001100010101010100101010110111010101001111011; end
            7'd49 : begin out <= 64'b0001101000000110101001011111100010101001100110110000111101011000; end
            7'd50 : begin out <= 64'b0010100011011010001000110100110000100100001000101010100110011001; end
            7'd51 : begin out <= 64'b1010101111110110101010000100101100101011001000011010010101001001; end
            7'd52 : begin out <= 64'b0010101111001101101011000110000110100100110101001010100001000110; end
            7'd53 : begin out <= 64'b0010100000110010101010001001100010100111111101111010101011111110; end
            7'd54 : begin out <= 64'b0010010011011110001001000000000110101001010111111010000101011011; end
            7'd55 : begin out <= 64'b0010011001000110100111110110011000100100011111111010100111011111; end
            7'd56 : begin out <= 64'b0001110010110011001010001101111100100101100101111010001001111111; end
            7'd57 : begin out <= 64'b0010100011100010001010110000001110100100100000110010011110100110; end
            7'd58 : begin out <= 64'b1001111100010001101010011001100110100111110000111010101110000100; end
            7'd59 : begin out <= 64'b0001101000000000101001000011111000101000100000100010000001101101; end
            7'd60 : begin out <= 64'b0001111101111011001001100010011100101000011011100010100001011100; end
            7'd61 : begin out <= 64'b1001110001000010001010100110111010101001001101000010001000110110; end
            7'd62 : begin out <= 64'b0010100001000101101000011111110100100110011110010010100011101110; end
            7'd63 : begin out <= 64'b0001110000001100001010111100011000100100101101001010001001100000; end
            7'd64 : begin out <= 64'b1010101011000011101010110001100100101001101101111010110001111000; end
            7'd65 : begin out <= 64'b1010101000111101001010100111011010101001010111000010101010101010; end
            7'd66 : begin out <= 64'b0001111010110101001010111011110100010110000001010010101111010011; end
            7'd67 : begin out <= 64'b1010000100101010101001011010100100101010110111100010100101001000; end
            7'd68 : begin out <= 64'b0010010100110111101010111101101010101000110111010010100001010011; end
            7'd69 : begin out <= 64'b0010011101001100001001100010000100101000101001010010101100110101; end
            7'd70 : begin out <= 64'b1010100110011010101001011111111100011111010011010010101010000000; end
            7'd71 : begin out <= 64'b1010101001101111001010001001110110101010010001010010101100100111; end
            7'd72 : begin out <= 64'b1010010111110011101001011111000100100101010111100010000001111001; end
            7'd73 : begin out <= 64'b0010100011101000101010010111110110100101110100001010011111100000; end
            7'd74 : begin out <= 64'b0010010011110000001001010011110110100111111000000010101100101010; end
            7'd75 : begin out <= 64'b1010100111100001101001101110111110101001001000001010011001110101; end
            7'd76 : begin out <= 64'b0010100111110000101011000111011100100000100001001010101010011011; end
            7'd77 : begin out <= 64'b1010100001011001001001111111111000100001110000010010011001001101; end
            7'd78 : begin out <= 64'b1010001001001101101010110100010010101011100011110001110101011010; end
            7'd79 : begin out <= 64'b1010100001110101101010001011100010100011100011010010101110001111; end
            7'd80 : begin out <= 64'b1010100000100001001010001000110010100001110100110010101110001111; end
            7'd81 : begin out <= 64'b1010101000101000001010000111101010100001111111111010001010011000; end
            7'd82 : begin out <= 64'b0010001010100010001000100110111000100101110100000010110000010001; end
            7'd83 : begin out <= 64'b0010100101101111001010000100100110101000001110100010011101110001; end
            7'd84 : begin out <= 64'b0010001001011111101010010111101010100101111110011001111001001111; end
            7'd85 : begin out <= 64'b0001011001000100101010100101111000100100100010001010011000000100; end
            7'd86 : begin out <= 64'b1010011110011100001010011101010000100110010110000010100110000001; end
            7'd87 : begin out <= 64'b0010100001001000101010011110011100101011101110101001110001100111; end
            7'd88 : begin out <= 64'b0001101110111101001010111011001010100101110001010010101100100111; end
            7'd89 : begin out <= 64'b0010100110110011001000001001001000100010110100000010001010110000; end
            7'd90 : begin out <= 64'b1010101111110110001010100011100010101001010000011010101110000111; end
            7'd91 : begin out <= 64'b1001011111011000001010001111111110101010001011110010010000001010; end
            7'd92 : begin out <= 64'b0010110000000010001000101001000010100011010101111010011001101010; end
            7'd93 : begin out <= 64'b0010010011111001100111001101111010101000010101110010101101111001; end
            7'd94 : begin out <= 64'b0010100110100100001001111000000000011110100011111010000110010100; end
            7'd95 : begin out <= 64'b0001110010100001001010000000110100101011101101100010000011010010; end
            7'd96 : begin out <= 64'b1010011010100001101000000000100100101011111001001010010100001110; end
            7'd97 : begin out <= 64'b0010000001010010100111101011001000101010101110111010101111110010; end
            7'd98 : begin out <= 64'b0010100001101001101000000111101100011011100111000010100000100100; end
            7'd99 : begin out <= 64'b0010011010010000001010001100000110101001010110011010011100111000; end
            7'd100 : begin out <= 64'b1010100111100001101010100001110000101000010010001010100110001101; end
            7'd101 : begin out <= 64'b1010100100110101101001101011010100101011000010110010010110101110; end
            7'd102 : begin out <= 64'b0010011101110111001001000111001010100101110110011010100011011001; end
            7'd103 : begin out <= 64'b0001111110101011101001100101101000101001110100001001100100100111; end
            7'd104 : begin out <= 64'b1010100010110101101010100100010110101001011001001010010011001111; end
            7'd105 : begin out <= 64'b1010000011011000101000110111111100100100011101011010010001100011; end
            7'd106 : begin out <= 64'b1010100011101110101010110111101100101011100001011010101000110010; end
            7'd107 : begin out <= 64'b1010100001101000001010011100100110101010100010101010011000000110; end
            7'd108 : begin out <= 64'b0010000010001000101011000111100110101000001001110010010100100000; end
            7'd109 : begin out <= 64'b1010100000011100001001001011011100100101011111000010100110000111; end
            7'd110 : begin out <= 64'b0010100001101000101010100000110000101001001000110010100111001010; end
            7'd111 : begin out <= 64'b0010010010001100001010001100011100101010101100001010101111001111; end
            7'd112 : begin out <= 64'b0010100011101100101010101111000110010111000001101001000101000011; end
            7'd113 : begin out <= 64'b0001110101111110001010110101001010101000001010101001011101100000; end
            7'd114 : begin out <= 64'b0010100011011010101000101110100110101010010011101001110000011001; end
            7'd115 : begin out <= 64'b0010010111101101001001001100111110101011000111010010011111010110; end
            7'd116 : begin out <= 64'b1010001110010111001010100000110100101011000000100001101000001111; end
            7'd117 : begin out <= 64'b1010100000110111101001100011111000101011000011100010010100110111; end
            7'd118 : begin out <= 64'b1001001110111100101001110001110010101001000100101010100101100000; end
            7'd119 : begin out <= 64'b0010010111110110001001001001101000101010001000111010001010011111; end
            7'd120 : begin out <= 64'b0010101000111001101010010110100010101001100011111010011001011010; end
            7'd121 : begin out <= 64'b1001100010000111001000010010111000101010010100100010101011100010; end
            7'd122 : begin out <= 64'b0010001101111001101001100111011100100100100100011010011001011000; end
            7'd123 : begin out <= 64'b0010101000111110001010011000001110101010110101010010000000011100; end
            7'd124 : begin out <= 64'b0010011101101000101010011010110000101001100100101001100110101011; end
            7'd125 : begin out <= 64'b1010101000000011001001000010001110100111111111101010011001010001; end
            7'd126 : begin out <= 64'b0010101100110000001000010101001100100110110011001010101000000100; end
            7'd127 : begin out <= 64'b1001010111010000001010110001000100011101110100000010001111001111; end
        endcase
    end
end
assign data = out;

endmodule //gemm3B
