
module gemm2B (
    input         clk,
    input         rst,
    input  [13:0] addr,
    output [63:0] data
);

reg [63:0] out;
always @(posedge clk or posedge rst) begin
    if (rst) begin
        out <= 0;
    end
    else begin
        case (addr)
            14'd0 : begin out <= 64'b1010100001011010101010011101010100101001010000110010101101001000; end
            14'd1 : begin out <= 64'b0001111110000111001010010011010000101010110110000010100110111001; end
            14'd2 : begin out <= 64'b0010001111001111001000001111110100100010100110000010101001111110; end
            14'd3 : begin out <= 64'b1010100110110010101010110110010000101000101011010010010001101000; end
            14'd4 : begin out <= 64'b1010010011001100101000011110011110100100111110010010101000101100; end
            14'd5 : begin out <= 64'b0010101000010100001000011011010000101011011010010010100000110000; end
            14'd6 : begin out <= 64'b1001110110000101101000100100001110101011110101101010001000101100; end
            14'd7 : begin out <= 64'b0010101110100111000110010110010000100010100101110010010011101001; end
            14'd8 : begin out <= 64'b0010100010011110101000011011100100011001000000111010100101111110; end
            14'd9 : begin out <= 64'b0010101001010010001001101111111100100100110101000010100111110000; end
            14'd10 : begin out <= 64'b0010001110110101101010101001110100101011011111000010011100110011; end
            14'd11 : begin out <= 64'b0010010101100010001010100100101010100001100100101010000110101111; end
            14'd12 : begin out <= 64'b1010101001110011101001010111110000100000001010100010100111000010; end
            14'd13 : begin out <= 64'b0010101001001010001010001010011100100110011000000010000010100100; end
            14'd14 : begin out <= 64'b0010010101110001101010010111100000101001111011000010010010011111; end
            14'd15 : begin out <= 64'b1010010011110000101010000110010000101000010111100001100101110010; end
            14'd16 : begin out <= 64'b1010101111001111001001110100000110011100010101000010011000000000; end
            14'd17 : begin out <= 64'b1010101111011001001001001100001000101010001011011010010010010111; end
            14'd18 : begin out <= 64'b0010100110100011101000011010101000101011000101110010010010110100; end
            14'd19 : begin out <= 64'b0010010011000001001001100101000010011100000101110001101110100001; end
            14'd20 : begin out <= 64'b1010101000001011100111110001011100101011011010101001010101100100; end
            14'd21 : begin out <= 64'b1010010010100111001010111111111010100111011001000010101011101110; end
            14'd22 : begin out <= 64'b1010001101101011001010100001101100100111110101111010101001010001; end
            14'd23 : begin out <= 64'b0010101100010101001001011101000110101010111011111010100111101111; end
            14'd24 : begin out <= 64'b0010000001111111101010100111000110011011001110010010010110110100; end
            14'd25 : begin out <= 64'b1010011101010110101001000001011110101010000010110010100010100010; end
            14'd26 : begin out <= 64'b0001111110010001001010010011101010100100010000111010011001101111; end
            14'd27 : begin out <= 64'b1010011010100001101001100000010000100011111010010001110001000010; end
            14'd28 : begin out <= 64'b1010101001010000101001100001101000101010100000000010011001110011; end
            14'd29 : begin out <= 64'b1010011001111100001001110000000000101001010110111010101010011001; end
            14'd30 : begin out <= 64'b0010011000100100101010010001101010101001110000011010100100011001; end
            14'd31 : begin out <= 64'b0010011100001111001001010001011110100101100100011010100010001110; end
            14'd32 : begin out <= 64'b0010101101000001000111111100100010101010010010110010110000010001; end
            14'd33 : begin out <= 64'b0010010101110011101001001000000000101011110011001010011101001111; end
            14'd34 : begin out <= 64'b0001111000001110101000111011111110101010001111011010000001001111; end
            14'd35 : begin out <= 64'b0010101100011101101000111001101110010100011011010010011011101101; end
            14'd36 : begin out <= 64'b0010010001001100100111000100010000101010010001010010100000101111; end
            14'd37 : begin out <= 64'b0010011001100111101010001001111000011011010100110001111010111000; end
            14'd38 : begin out <= 64'b1010101011110011101001010100110100100100001010100001111111010001; end
            14'd39 : begin out <= 64'b1010101101001110001001111111100010101001101000101010100010101000; end
            14'd40 : begin out <= 64'b1010101011101111101010111001000110100100001111110010000111010100; end
            14'd41 : begin out <= 64'b1010101110010001101001101111101110100010110011011010101001101101; end
            14'd42 : begin out <= 64'b1001101011101011101010111101110000011100110100101010010100100000; end
            14'd43 : begin out <= 64'b1001011010001001101010100100100010100001010101101010010110100010; end
            14'd44 : begin out <= 64'b1010101001111100101001101011010010100001100111101010010010100000; end
            14'd45 : begin out <= 64'b1010010010110010100000000000111100101000100111100010000011000001; end
            14'd46 : begin out <= 64'b0010101100011110101010100111111000100110100110100010100011101001; end
            14'd47 : begin out <= 64'b1001110100011110101010111111000100100001000010101010010101100011; end
            14'd48 : begin out <= 64'b0010101101111000001010101100011010100010111101101010110000010000; end
            14'd49 : begin out <= 64'b1010011001010011101000011111000100101001110111100010100011100001; end
            14'd50 : begin out <= 64'b1010101011000001100110010011100010101000110100010010101100110001; end
            14'd51 : begin out <= 64'b0010100010111110101010111001001010101010000110101010011000001011; end
            14'd52 : begin out <= 64'b0010101101010100001001000010000000101000101110110010011100011111; end
            14'd53 : begin out <= 64'b0010101010011000101010010100011010101001111011000001011001111110; end
            14'd54 : begin out <= 64'b0001111100011111101001000010100010101011101011011010100010011001; end
            14'd55 : begin out <= 64'b1010100010100101001001011011011000101001100110000010101101100001; end
            14'd56 : begin out <= 64'b0010011101101000101010100010111000101011001010100010100101000111; end
            14'd57 : begin out <= 64'b1010100110111011101010111011000010101010001100100010101110011011; end
            14'd58 : begin out <= 64'b0010101000000011101001010010011110100000111110000010101111110011; end
            14'd59 : begin out <= 64'b1010101011111111001010010010000010101010000010111010100111001010; end
            14'd60 : begin out <= 64'b0010001100111110101001000111110110100011001111111010001010110011; end
            14'd61 : begin out <= 64'b1010100111110111001001100110010010100110011111001001110110011000; end
            14'd62 : begin out <= 64'b1001111010001100101010010000010110010110001100010010101110110001; end
            14'd63 : begin out <= 64'b1010101100011111101001001010110010101011111100100010010001100010; end
            14'd64 : begin out <= 64'b0010100001010111101010100111100110101000110110101010100011100111; end
            14'd65 : begin out <= 64'b1010101000010101001010101010110010101011101000001010011001011111; end
            14'd66 : begin out <= 64'b0010101000011101101001111110011000101011010011000010010100100110; end
            14'd67 : begin out <= 64'b1010000110010101101001110011101010101000110010000010100010010010; end
            14'd68 : begin out <= 64'b1001100001001101101010110100101100101000001110010010100000000110; end
            14'd69 : begin out <= 64'b1001110010100010001010000101100100100110011100001010100110111111; end
            14'd70 : begin out <= 64'b1010010001011111001001101100011010101011110101001010101111000111; end
            14'd71 : begin out <= 64'b1010010000110100001010101100001100100100100000011010101101001011; end
            14'd72 : begin out <= 64'b1010011011111000101010001010011000101010110010001010011001001101; end
            14'd73 : begin out <= 64'b0010100111001111001010001101000010101000001010001010101001001100; end
            14'd74 : begin out <= 64'b0010010011011101001010000010100000101001101111101010010001110100; end
            14'd75 : begin out <= 64'b1010101000111001001000110111000010101010001111101010001110011101; end
            14'd76 : begin out <= 64'b0010000110001111101000000101110100101001001111011001100111100010; end
            14'd77 : begin out <= 64'b1010011011010010101010000001010110101001011011110010101011011110; end
            14'd78 : begin out <= 64'b1010101100101000100111000001010010011101100110000001111110101001; end
            14'd79 : begin out <= 64'b1010101010100100101001100001010010100010111100001010011010111111; end
            14'd80 : begin out <= 64'b0001110101110110000100011011100000101001101100101010100000100000; end
            14'd81 : begin out <= 64'b1010010010011110101000010100110110010100010100111010011000100010; end
            14'd82 : begin out <= 64'b1010010000111000101010101000001000101010000000111010010000001000; end
            14'd83 : begin out <= 64'b0010101000011001001010011110111110100101010001001010011011000101; end
            14'd84 : begin out <= 64'b1010100001110101001000110011011100100000000011011010100110110011; end
            14'd85 : begin out <= 64'b1010100011011100100110101100000010101000100011111010101111101001; end
            14'd86 : begin out <= 64'b0010000101110111001010101101101110100000001011000010100111000100; end
            14'd87 : begin out <= 64'b1010100100011010000110001110110110101010111101011010011000110001; end
            14'd88 : begin out <= 64'b0010000001101001101001010001101110100100101110001010010100000110; end
            14'd89 : begin out <= 64'b1001110000011001001010000111100010100110011011111010011011101110; end
            14'd90 : begin out <= 64'b0010001101100111001000011110110110101000001001001010100100000100; end
            14'd91 : begin out <= 64'b0010001011010111001001101110000010100101110101100010011100001100; end
            14'd92 : begin out <= 64'b1010101011101111001010100000101000100111000000101010001000000100; end
            14'd93 : begin out <= 64'b1010100000011101101010101000010010101000111000111010011100100010; end
            14'd94 : begin out <= 64'b1010101000001110001010111010111100101000111010011010101011010011; end
            14'd95 : begin out <= 64'b1010011011010101100111000000110010101011101010001010101010011000; end
            14'd96 : begin out <= 64'b1010001101110011000111000001010100100100111101010010011011011110; end
            14'd97 : begin out <= 64'b0010100101101000101001001010100110101011100011001010101000100001; end
            14'd98 : begin out <= 64'b0010100111010110001001001001000000010110111000111001100101101100; end
            14'd99 : begin out <= 64'b0010011110001010001010010011000000100100111111011010010100001111; end
            14'd100 : begin out <= 64'b1010101010001111001010011000111010101000010000001010101111100111; end
            14'd101 : begin out <= 64'b1010101110001111101010000010001010100110110100001010101010100101; end
            14'd102 : begin out <= 64'b0010100111111001101010001101000100101011001110110010011010010010; end
            14'd103 : begin out <= 64'b1010100011111101001010011110011000101000011101100010000100101110; end
            14'd104 : begin out <= 64'b0001111001101010101010000101100000101011111100000010011100011110; end
            14'd105 : begin out <= 64'b1010101011100011001010001000001010101001010110001001110000001000; end
            14'd106 : begin out <= 64'b0001100111101110101001011111001010100111011011001010100100100111; end
            14'd107 : begin out <= 64'b1010001101000001001001001110111100101010000001100010011000100000; end
            14'd108 : begin out <= 64'b1000100001101111101010000100110010011001101011010010101001011000; end
            14'd109 : begin out <= 64'b0001001000110110101000011100101100101011010100100010011011010100; end
            14'd110 : begin out <= 64'b1010101100011100001001101101111110101010101101100010101001101011; end
            14'd111 : begin out <= 64'b1010010101110011001000011010111010101010100011100010010011100100; end
            14'd112 : begin out <= 64'b1010101101010000101010000111011000101001110001101010100101000100; end
            14'd113 : begin out <= 64'b1010010100000001001001001000100100101000100001111010100111000110; end
            14'd114 : begin out <= 64'b0010101110111000101010110000101110100011011111111010100010001110; end
            14'd115 : begin out <= 64'b0010101111001001001010010110010100101001100110100010100101001000; end
            14'd116 : begin out <= 64'b1010000001111000001010111101101110101001000111101010101100010110; end
            14'd117 : begin out <= 64'b0010100101000110001010011001000110100110100100000001110000111100; end
            14'd118 : begin out <= 64'b0010010110000011001001111001010110101010110011000010101111110100; end
            14'd119 : begin out <= 64'b1010100011001110001001101111111110100100100010110001110010111111; end
            14'd120 : begin out <= 64'b0010100010100110101001001100011100101001110110101010101011110000; end
            14'd121 : begin out <= 64'b1010010000001011100110101111000010101011111001100010101010111110; end
            14'd122 : begin out <= 64'b1001100000010010101010101110010000101011001101100010011110101100; end
            14'd123 : begin out <= 64'b1010001000111000101001010011011010101000100001111010010001000011; end
            14'd124 : begin out <= 64'b0010100011111001001010100111001010010110000001100010101001001000; end
            14'd125 : begin out <= 64'b1010100111010110001010100000100000101000110101001010000011111110; end
            14'd126 : begin out <= 64'b0010010011011001100110100001100100100111011010110010000101100011; end
            14'd127 : begin out <= 64'b1010100110011101001001111101001010011101110101000010101111010011; end
            14'd128 : begin out <= 64'b0010100101011111101010000110011100100000100011010010011001001001; end
            14'd129 : begin out <= 64'b0001011110010001001010011111001010100101010111010010011101010000; end
            14'd130 : begin out <= 64'b1001011000110110101010001010111110100101000111000010100011011010; end
            14'd131 : begin out <= 64'b1010010010000101100110110110000100101011000101011010010101100011; end
            14'd132 : begin out <= 64'b0010100001101101100110010001010100100011111101010010101110101011; end
            14'd133 : begin out <= 64'b1010011011000111001001100101011100100101011000000010011111011101; end
            14'd134 : begin out <= 64'b1010000101011001101001111101010100100111011100011010000110010011; end
            14'd135 : begin out <= 64'b1010100000100001101001010011000000101011000010011010101110010110; end
            14'd136 : begin out <= 64'b0010100111111000001010001010101010100110000111010010101011001110; end
            14'd137 : begin out <= 64'b0001110010111011101000100111001000101000111010101010001011000011; end
            14'd138 : begin out <= 64'b1010011001110011001001010001011100100100001111000010101100000111; end
            14'd139 : begin out <= 64'b0010101100111110101010101010001010100001101111001010010100010001; end
            14'd140 : begin out <= 64'b1010001110000011001000000010111110100111100110101010100000011001; end
            14'd141 : begin out <= 64'b1010000001010001001010111010000100101010101100011010011011110110; end
            14'd142 : begin out <= 64'b0010010111010110001010100001110010101010011011101010101011011010; end
            14'd143 : begin out <= 64'b1010000001111001000110011010111100100010110000010010100110101110; end
            14'd144 : begin out <= 64'b1010101100100110101010111110000110100110111101100010100000110101; end
            14'd145 : begin out <= 64'b0010100110110110001010110011010100100100000111110010010000101111; end
            14'd146 : begin out <= 64'b0010100101001000001010110110111100101000100101001010101100010101; end
            14'd147 : begin out <= 64'b0001101001110010101000111101110010011110011111111010001011101000; end
            14'd148 : begin out <= 64'b1010000000111010001010111100011100100111010001101010100010101011; end
            14'd149 : begin out <= 64'b0010011011011110101010101110100000101000010111101010000000000010; end
            14'd150 : begin out <= 64'b0010101110011111001001111101100000101001101011110010100001010000; end
            14'd151 : begin out <= 64'b1010000100011100101001000110110010101000010101000010100100101101; end
            14'd152 : begin out <= 64'b0010000100101111001010011011100010100110000110101010100110100000; end
            14'd153 : begin out <= 64'b0010011111001000001010011101010010100001000000111010000011100010; end
            14'd154 : begin out <= 64'b1010100110000111101000011101111100101001111101011010101000111100; end
            14'd155 : begin out <= 64'b1010011100110101101001010010001010011100000000110010101100001011; end
            14'd156 : begin out <= 64'b0010100011110001101010000000001010101011111101101010001000110000; end
            14'd157 : begin out <= 64'b0010001001111001101010101010110100100110000001011010011001011111; end
            14'd158 : begin out <= 64'b0010100001101000001000001110100100100000001101111010101011101011; end
            14'd159 : begin out <= 64'b1010001110110110101010000001010000101001010111101010100101111001; end
            14'd160 : begin out <= 64'b0010000100100110101000000111010100100101001100000010101100011101; end
            14'd161 : begin out <= 64'b1010100100000101000100100011000000100101101010000010011000110000; end
            14'd162 : begin out <= 64'b0010101111000000101010110001010000010111101000011010001000111101; end
            14'd163 : begin out <= 64'b0001110110111001001001100011111110101001110110111010010011000000; end
            14'd164 : begin out <= 64'b1010100000111111001010000111111000100110100000100010100110000110; end
            14'd165 : begin out <= 64'b1010101001000010101010111100111100101001101100001010010010100110; end
            14'd166 : begin out <= 64'b1010100011011010001001111000111000101000001011000010101101000110; end
            14'd167 : begin out <= 64'b1010011011101111101010001100010000100111101011110010010001010101; end
            14'd168 : begin out <= 64'b1010100110101001001010000001010010100100000110110010011101000101; end
            14'd169 : begin out <= 64'b1010100100011001001010000010000010100100101110101010010101000100; end
            14'd170 : begin out <= 64'b0010011111100000001001101111101000101001001101110010101101100101; end
            14'd171 : begin out <= 64'b1010001100100110001010100010001010100111011000111001111000111010; end
            14'd172 : begin out <= 64'b1010011110000101101010101111101000011101010111010010101100001100; end
            14'd173 : begin out <= 64'b0010001000110111001010100100011000101000010111101010010000001111; end
            14'd174 : begin out <= 64'b0010100111011010100111011011111100101010010001011010101011111100; end
            14'd175 : begin out <= 64'b0010101111100010101001110100110100101000100111001001110001101010; end
            14'd176 : begin out <= 64'b0010000100011000101010011000010000101000000101001010010111010001; end
            14'd177 : begin out <= 64'b0010011001011011000110100001010010100011001000100010101001111111; end
            14'd178 : begin out <= 64'b0010101001111110001000010101100110101010001000101010101001101101; end
            14'd179 : begin out <= 64'b0010101011110101101010111010101000011100101010011010101001111100; end
            14'd180 : begin out <= 64'b1010101100111110001001001011101010100100110100000010100010110100; end
            14'd181 : begin out <= 64'b0010101101000100000101110011001000000001101101011010100110110110; end
            14'd182 : begin out <= 64'b0010011011100101101001000100110000101001011001110010010011111011; end
            14'd183 : begin out <= 64'b0010011111010011101010111101101010011000101100111010100111110100; end
            14'd184 : begin out <= 64'b1010100001001110101001000011000010101001011101101010100110110011; end
            14'd185 : begin out <= 64'b0010001101101001001010111100110010101000111000101010101000010011; end
            14'd186 : begin out <= 64'b0010000010100001001000111101111100101001110101111010110000000000; end
            14'd187 : begin out <= 64'b1001010001100111001010100000000100101000111101000010100110000111; end
            14'd188 : begin out <= 64'b0010101010110101101010011100000010100111100010110010100101111111; end
            14'd189 : begin out <= 64'b1010100000010110101010010111101110101011111111100010100000010111; end
            14'd190 : begin out <= 64'b1010011111110001101010000100110010011110001101110010010110110100; end
            14'd191 : begin out <= 64'b1010101010011010001001010111011100100110000111011001110011001100; end
            14'd192 : begin out <= 64'b1010101000100111101000100110110000100100111100010001011010010000; end
            14'd193 : begin out <= 64'b1010100100011000001010110110001110001011111011111010100010011100; end
            14'd194 : begin out <= 64'b0010101100100100101010001100110010010010111111110010101010110000; end
            14'd195 : begin out <= 64'b0010100100010110001010111111001100100101000011001010010111010001; end
            14'd196 : begin out <= 64'b1010010110100111001010101100111010101000110110010010100010011110; end
            14'd197 : begin out <= 64'b1010101100010111101001100111011010100110000111101001101001000011; end
            14'd198 : begin out <= 64'b1010101101110011001001101100011010101001101110110010011001101001; end
            14'd199 : begin out <= 64'b1010100010101100101001000011111000101011110100110010001001001101; end
            14'd200 : begin out <= 64'b0010011100100000000101010111101010100111000100101010101001111000; end
            14'd201 : begin out <= 64'b0010010010101000001010111001111000101001011110100010101011110110; end
            14'd202 : begin out <= 64'b0001111000010010101010111111010100100111011101111010100101000001; end
            14'd203 : begin out <= 64'b0001100010111110101010101011001000101011111011000010011100100011; end
            14'd204 : begin out <= 64'b0001101101100010001001101110000100101011010100010010100011110000; end
            14'd205 : begin out <= 64'b1010010100001010001000011010101100101000000010010010100011111000; end
            14'd206 : begin out <= 64'b1001111110000100101001111111011100101010001001111010011110001111; end
            14'd207 : begin out <= 64'b1010101100100001000101101000011110101001011100100010011110100100; end
            14'd208 : begin out <= 64'b1010010010111101001001001001100010101001101000000010101000011101; end
            14'd209 : begin out <= 64'b0001100011111000001010001001001000100110100100010010101001100111; end
            14'd210 : begin out <= 64'b0001000010000111001010000011010000101000110000100010000011111100; end
            14'd211 : begin out <= 64'b1010101000011010101010100010110000100001010101000010000101000100; end
            14'd212 : begin out <= 64'b0001101100111110100100010011110010010001100010011010100111011000; end
            14'd213 : begin out <= 64'b1010100101110110001010110001101100011111100000001001111110010111; end
            14'd214 : begin out <= 64'b0010011000001110001010111110011100100100010001101010100010101100; end
            14'd215 : begin out <= 64'b1010010100111110001001001001010110100101011111011010010110111100; end
            14'd216 : begin out <= 64'b1010011011001000001001111010100000100001110110000001010010010010; end
            14'd217 : begin out <= 64'b1001110010101111001000110100010000101011110100101010000100011000; end
            14'd218 : begin out <= 64'b0010101110011111001010110011101100011100000001110010010011010101; end
            14'd219 : begin out <= 64'b1010011111100101100111100101110000101010110110011010010101100110; end
            14'd220 : begin out <= 64'b1001110011001011001010010001100000101001001011110010011101010010; end
            14'd221 : begin out <= 64'b1010011000001000101001001100111010011001100010110010101010100011; end
            14'd222 : begin out <= 64'b1010101011110111000011110010101000101001000010010010100100100010; end
            14'd223 : begin out <= 64'b0010101011010001101000100000010000101001010110010010001110101001; end
            14'd224 : begin out <= 64'b1010100010001110001001111001110110101010111000101010011111011010; end
            14'd225 : begin out <= 64'b1001100111101100100100111000111100101011001011110010000100110001; end
            14'd226 : begin out <= 64'b1010011110111100000111011110111100101010001101000010011111000001; end
            14'd227 : begin out <= 64'b0010100110011001001010110001100110011011100110111010101011001000; end
            14'd228 : begin out <= 64'b0001100101111100001001110101010110101011001001001010000101001001; end
            14'd229 : begin out <= 64'b0010100110001000101001110010100100101000001100000010101011011001; end
            14'd230 : begin out <= 64'b0000111010111001101010110010011010101010101101110010100110011010; end
            14'd231 : begin out <= 64'b0010010000101110000110100111011100101000101000010010001000010010; end
            14'd232 : begin out <= 64'b0010100010110100001001111010010000101010010111001010101110000100; end
            14'd233 : begin out <= 64'b1010101011010011001010010101011000100000100001100010001101100100; end
            14'd234 : begin out <= 64'b0010101000001001101010111011010000101010100110101001110001010011; end
            14'd235 : begin out <= 64'b1010100101111100101010100000001100101000000011011010101010110011; end
            14'd236 : begin out <= 64'b0010101111110001101001010001010010101011101111010010010001101111; end
            14'd237 : begin out <= 64'b1010101101100110001010101101001110100111011001111001101011111010; end
            14'd238 : begin out <= 64'b0010011011001000101010010001100100101011011111100010010000010000; end
            14'd239 : begin out <= 64'b1010001011110100100101100110000010100111100101101010101101101000; end
            14'd240 : begin out <= 64'b1001111110111110101010010010101110100110110010110010100011110000; end
            14'd241 : begin out <= 64'b0010011000100111100111010010010000100100010110111010101000011100; end
            14'd242 : begin out <= 64'b0010010100110111001000010111100110101000100101011010101010010000; end
            14'd243 : begin out <= 64'b1010001101001101001001100000110100100110100011101010101110110110; end
            14'd244 : begin out <= 64'b0010100111011100001010001100010010011000110000100010001001000001; end
            14'd245 : begin out <= 64'b0010101011101100001010101011101010100101010101101010010111010110; end
            14'd246 : begin out <= 64'b0010101100110010000110111011100000101011001011111010101100111010; end
            14'd247 : begin out <= 64'b0010101000001011100111101110010000101001110000111010101000111111; end
            14'd248 : begin out <= 64'b0010101110001101001010001110010100010100011110101010001001000001; end
            14'd249 : begin out <= 64'b1001111100111011100111011000100110101000101001110010101001001011; end
            14'd250 : begin out <= 64'b1010101110100111001001000101111100101011011011010010010110110111; end
            14'd251 : begin out <= 64'b1010101100101010101001001101111110101010000011110010101110011101; end
            14'd252 : begin out <= 64'b1010100001001111000111010100101100101000101011101010101000110111; end
            14'd253 : begin out <= 64'b0010000001011101001010010001001100101000111010101010101010001101; end
            14'd254 : begin out <= 64'b1010100110110111001010010101101100101000100101010010100011111011; end
            14'd255 : begin out <= 64'b1010101000111001001000110111111000101001001011001010000101100111; end
            14'd256 : begin out <= 64'b0010011100010000001001010011000110101011000011100010010111000001; end
            14'd257 : begin out <= 64'b0010100100101011101000010000000000101011111101000010101011111010; end
            14'd258 : begin out <= 64'b0010101101001111101010011011111110101011100100010010100010101011; end
            14'd259 : begin out <= 64'b1010100001101110101010010011100110101010010100101010100001010011; end
            14'd260 : begin out <= 64'b0010100110101110101000100011101110101011110100011001111100101100; end
            14'd261 : begin out <= 64'b0010000100001000001010001010000010101010111100000010100111100110; end
            14'd262 : begin out <= 64'b1010101011110110001010110000101100101001110011001010010100000000; end
            14'd263 : begin out <= 64'b0010001110000000001010010000010110101010011011011010100010001111; end
            14'd264 : begin out <= 64'b1010010100110011001010110001100100101000010110010001110010100100; end
            14'd265 : begin out <= 64'b0000111110110111101010001011000000100100110111111010100010110101; end
            14'd266 : begin out <= 64'b1010001011001001101010010001110100011001101011111010101110111001; end
            14'd267 : begin out <= 64'b1001110011111000101010001011001000101000011010011010101011000100; end
            14'd268 : begin out <= 64'b0001100001011001001001110111011100101010100110011010001011010001; end
            14'd269 : begin out <= 64'b0010100000000101101010001001000000101001100011000010100010110000; end
            14'd270 : begin out <= 64'b1010010100101000000100000001011010101010010111000010100010110110; end
            14'd271 : begin out <= 64'b1010100001101010001000100110000010101011100111101010010010011101; end
            14'd272 : begin out <= 64'b1010001101111110001010110011101100101011011001010010100001010111; end
            14'd273 : begin out <= 64'b1010011110101001001001010101101000101011100001111010010000101000; end
            14'd274 : begin out <= 64'b0010010101000111001000010111001010101001011001111010000101110000; end
            14'd275 : begin out <= 64'b1010010000010000001010000100100010101000001110000001000100110010; end
            14'd276 : begin out <= 64'b0001101000111110101000110110010100101000110000011010101111101000; end
            14'd277 : begin out <= 64'b0000000101100011101010111010010010100010111010101010100100010110; end
            14'd278 : begin out <= 64'b0010010110110001001010111110010000101010000110101010100011101111; end
            14'd279 : begin out <= 64'b0010101101011001101001011011111100101001110010111010101001011000; end
            14'd280 : begin out <= 64'b1010100111011010101010010011010010101000001000110001000111111001; end
            14'd281 : begin out <= 64'b0010011111001010001000111111010010101010100111010010101110010011; end
            14'd282 : begin out <= 64'b1010101100111000000110010101110110101001000011100010101111010010; end
            14'd283 : begin out <= 64'b0010011110000001000110110111010000101010011100101010101100001110; end
            14'd284 : begin out <= 64'b1010101011110111101010111101100010100010110000000010101111010000; end
            14'd285 : begin out <= 64'b0001100101001000101001011000100010100111111000101001101100000110; end
            14'd286 : begin out <= 64'b0010101110000000001010001110111100101010100101111010001110010101; end
            14'd287 : begin out <= 64'b1010010010110111001001100010101010100111101000011010000111001101; end
            14'd288 : begin out <= 64'b1001110111111001001000000000111010101011100010011001101011010010; end
            14'd289 : begin out <= 64'b1010100110011100001010011100001100101010110001100010000000010010; end
            14'd290 : begin out <= 64'b1001111010010010101010010001110010100100000100111010011001000100; end
            14'd291 : begin out <= 64'b0010110000111010001011000101100000101001111110110010100001010100; end
            14'd292 : begin out <= 64'b1010101000011111001010010000100000101010001001001010100001101001; end
            14'd293 : begin out <= 64'b1010101111111001001001111101011000101011000110111010011111011001; end
            14'd294 : begin out <= 64'b1010000110111100001001110100101110101000100100100010010000100110; end
            14'd295 : begin out <= 64'b1010001001101101101010101111011110101001111001110010100010011111; end
            14'd296 : begin out <= 64'b0001011100110001001010001001010000101011110000010010001110111110; end
            14'd297 : begin out <= 64'b1010101100101111101010010100000000100110111011101010100100100010; end
            14'd298 : begin out <= 64'b0010100110111100101010110101011010100110100100100010010100110001; end
            14'd299 : begin out <= 64'b0001010100011011001010100101111010011100111100010010100111110011; end
            14'd300 : begin out <= 64'b0010101001110111101001110000000110101010001100110010100010011111; end
            14'd301 : begin out <= 64'b1010011111100111101001011000010110101001000000011010100001111111; end
            14'd302 : begin out <= 64'b0010011000100010000111100111001110010101011111011010001000001100; end
            14'd303 : begin out <= 64'b0010001110110000001010111011111000101001001010001010010101011101; end
            14'd304 : begin out <= 64'b0010010001011100101001011010000110100010101111010001100110100101; end
            14'd305 : begin out <= 64'b1010010001011110101001110100111100100101101110110010100010111001; end
            14'd306 : begin out <= 64'b1010100000101100001000100011101010101011010111000010101100110101; end
            14'd307 : begin out <= 64'b1010101111110111101001101101010000101001100001101001101001101011; end
            14'd308 : begin out <= 64'b1010100000110100001010101001001100010110111100010001111001010010; end
            14'd309 : begin out <= 64'b0010011101101010001010011111000100100110000110100010100100100111; end
            14'd310 : begin out <= 64'b0010010011011001001010010110001010011100100100111010100100000111; end
            14'd311 : begin out <= 64'b1010101011111001101000001000100100100100001111111010001001000111; end
            14'd312 : begin out <= 64'b1010001100111011101001101110010010101001110001011010100011000000; end
            14'd313 : begin out <= 64'b1010011110011100100111010101110000101000010010011001101101110110; end
            14'd314 : begin out <= 64'b1010100011111101101010100000010000100110000101101010010111101000; end
            14'd315 : begin out <= 64'b1010011001010001101001100101101110100100010100110010101100001101; end
            14'd316 : begin out <= 64'b1010010110100101101010110110100110101010100100100010000010100001; end
            14'd317 : begin out <= 64'b1001110011000110001010011001010010101001110011010001110110001111; end
            14'd318 : begin out <= 64'b1010101100000011001000101100111000101000100011000001101110101111; end
            14'd319 : begin out <= 64'b1010011110111011101010011011111000100010110011000010000011000011; end
            14'd320 : begin out <= 64'b0010101111011000100111001110100000101010010101101010101110111110; end
            14'd321 : begin out <= 64'b0010000010000011001001010101001110101010110001010010000100001010; end
            14'd322 : begin out <= 64'b0010101101011001001010110100111010000111010011011010101100000111; end
            14'd323 : begin out <= 64'b1010100001110000001010100100110010101001110000010010011000100110; end
            14'd324 : begin out <= 64'b1001110111111000101001111001111000101011011001100010100000100110; end
            14'd325 : begin out <= 64'b0001011010011111101010111110001100100111110010101010011011100010; end
            14'd326 : begin out <= 64'b0010101011010101001010011110011100101011011001001010001110001100; end
            14'd327 : begin out <= 64'b1010101101011101001001011010000010101001000001101010001001010110; end
            14'd328 : begin out <= 64'b0001111000101110101010001011101100100111100011001010001110100000; end
            14'd329 : begin out <= 64'b1010000110100110001010100100110100100011100001101010011100000010; end
            14'd330 : begin out <= 64'b0010101100110011101010001011001000100101110001101001101000101111; end
            14'd331 : begin out <= 64'b0010101101001010101010010010101100101000001011111010101110100110; end
            14'd332 : begin out <= 64'b0010100010001110101010000111011010101011110011010010100101100000; end
            14'd333 : begin out <= 64'b1001101000010010101000010011110010100000011010100010001011101111; end
            14'd334 : begin out <= 64'b1010001111010101001001000100010110101011000000100010100011110110; end
            14'd335 : begin out <= 64'b1010000011011101001010100011011010101001001101100010011010101101; end
            14'd336 : begin out <= 64'b0010100100100000101010100110001110100110100110101010101111011101; end
            14'd337 : begin out <= 64'b1000101011101000101010101110001000101011001001110001110011000110; end
            14'd338 : begin out <= 64'b0010100010100100000111101001111000101011101101000010100001111100; end
            14'd339 : begin out <= 64'b1010000000101001001001110010010010101001111100001001101110011101; end
            14'd340 : begin out <= 64'b0010101000111011001001110010011100100111110101000010101001101111; end
            14'd341 : begin out <= 64'b0010000001100101001010111001100100101001000100001010100110000110; end
            14'd342 : begin out <= 64'b1001110111111101001001100001010100011001100111100010100010000111; end
            14'd343 : begin out <= 64'b1010010010110110101010011100101110101001000100001010100100101001; end
            14'd344 : begin out <= 64'b1010100111000110000110111110101010101000001010010010101000010001; end
            14'd345 : begin out <= 64'b0010010111100010001001000001001100100101010011001010101010000011; end
            14'd346 : begin out <= 64'b0010011110101110001001101001000100101010101010101010000011110110; end
            14'd347 : begin out <= 64'b0010101010110101001010101101100100010100100101101010011111110110; end
            14'd348 : begin out <= 64'b0010011001000010100111010110000010101001100000101010100001001111; end
            14'd349 : begin out <= 64'b0010100000100110101010010111011000101001011110000010000111000110; end
            14'd350 : begin out <= 64'b1010010101110110101010110000001000101001001101110001010001100001; end
            14'd351 : begin out <= 64'b1010100100000110101011000110010110101000101110010010101000100001; end
            14'd352 : begin out <= 64'b1010010010110000101010011111010000010111011100000010100101000000; end
            14'd353 : begin out <= 64'b0001110110010110101001010100010000100000111100011010101000101000; end
            14'd354 : begin out <= 64'b1010010011100100001010011100111110101000100100001010101010011101; end
            14'd355 : begin out <= 64'b0010011000011100001010000001110110100111100011000010000001100101; end
            14'd356 : begin out <= 64'b0010000001000011101010011010111000100100010111000010101100100111; end
            14'd357 : begin out <= 64'b1010101101111100001010001111011000101010010101001010100100000101; end
            14'd358 : begin out <= 64'b1010100111110101101010001100100110010111000001101010010011010011; end
            14'd359 : begin out <= 64'b0010011001000101001010101000001000101001110000011010000001001101; end
            14'd360 : begin out <= 64'b1010011111111110001001101100011010011000111111000001111001101101; end
            14'd361 : begin out <= 64'b1001111001000110001000000101011110101011110001101010100000111010; end
            14'd362 : begin out <= 64'b0010010001011111000101000010011010100110110111111010100010111110; end
            14'd363 : begin out <= 64'b1010101000111100001010101011110100011100101100000010101001100110; end
            14'd364 : begin out <= 64'b0001110100010101001010011101010110101011111011100010100011101110; end
            14'd365 : begin out <= 64'b0010100111110101001010011101111110101010010011101010101000001111; end
            14'd366 : begin out <= 64'b1010100010011100000100001111110100100001101100011010000101100000; end
            14'd367 : begin out <= 64'b1001011101000100001000100110001000101010111100110010010010000010; end
            14'd368 : begin out <= 64'b0010101011101101101000000110010110101000110111101010101010000010; end
            14'd369 : begin out <= 64'b1010010010010110101010101100001110100100111011111010101011110011; end
            14'd370 : begin out <= 64'b0010000111101011001010101011010110101010000010101010101001010111; end
            14'd371 : begin out <= 64'b0010010001010010101000010101101100101011010100000010101111000000; end
            14'd372 : begin out <= 64'b1010101100110000101010110110010110101001001110111010011111110010; end
            14'd373 : begin out <= 64'b0010100001000111101000100011100110010111001101011010001101001010; end
            14'd374 : begin out <= 64'b1010101100010100101010111110001010100111110100011010100101111011; end
            14'd375 : begin out <= 64'b0010101110100100001010111011011000100011000100110010100100011111; end
            14'd376 : begin out <= 64'b0010100000011000101001110111110010101000010101100010011000001101; end
            14'd377 : begin out <= 64'b1010100010101001101010100001001000101011100011111010100011001101; end
            14'd378 : begin out <= 64'b0010101100000100101001000111010100101001000100111010011111101010; end
            14'd379 : begin out <= 64'b1010100111100111101010011010010110100100111111000010101111010110; end
            14'd380 : begin out <= 64'b1010101100101010101010100001101100011100011111110010100111001101; end
            14'd381 : begin out <= 64'b1010010110000110101001110001011000100110111101100010011101100101; end
            14'd382 : begin out <= 64'b0010011111001111100110101000111000101000110111110001011110011001; end
            14'd383 : begin out <= 64'b0010101000010011001000000100010100101001110101101010010100111110; end
            14'd384 : begin out <= 64'b1010100110111010100110010001001000101000001100111010101111001010; end
            14'd385 : begin out <= 64'b1010100100110110101010011110111110100101000100011001111111110101; end
            14'd386 : begin out <= 64'b1010011011101001100111110011110010101011010101100010101101100011; end
            14'd387 : begin out <= 64'b0010110001010010001010111111010100100001011110110010100100011010; end
            14'd388 : begin out <= 64'b1001111010010000101010000011011000011010010000111010101110111011; end
            14'd389 : begin out <= 64'b1010101001001111100111000111111010100011111101001010100100100101; end
            14'd390 : begin out <= 64'b1010100101110010101000001001100000100011111011010010101110100000; end
            14'd391 : begin out <= 64'b0001110110001001001001011000110010101011011011100010100111111000; end
            14'd392 : begin out <= 64'b0010100101010110001001111101010110101010010001100010100101100011; end
            14'd393 : begin out <= 64'b1010011011110000001010111111011100101000010000101010001000111001; end
            14'd394 : begin out <= 64'b1010011101111100101001010111111000101001101010100010000110111111; end
            14'd395 : begin out <= 64'b1010101111110100101010110110100110011110111110110010100000101111; end
            14'd396 : begin out <= 64'b0010001111001110001010000001001000100100000111110010101000000110; end
            14'd397 : begin out <= 64'b0010000011100010001001101101100110100100100110111010000111000011; end
            14'd398 : begin out <= 64'b1010100001011000001001000111000000101001001111011010000110000000; end
            14'd399 : begin out <= 64'b1010101011011110100111011101110110100001000111101001100110000010; end
            14'd400 : begin out <= 64'b1001101111011111101010000100110100100110010101111000111011100111; end
            14'd401 : begin out <= 64'b0010101011101001101010111101101110101001001111111010101101111000; end
            14'd402 : begin out <= 64'b0010101001010110101001100000010110100110010001110010100010101010; end
            14'd403 : begin out <= 64'b1001110000011111000101111111101010101010100010100010011010110000; end
            14'd404 : begin out <= 64'b1010010010000101101010101000010010101000011111001010001000000111; end
            14'd405 : begin out <= 64'b1010000111010010001000011001001110100000011010010001100101011001; end
            14'd406 : begin out <= 64'b1010011100001001101010000011000110011110110111001010000111000101; end
            14'd407 : begin out <= 64'b1010010001010001001000101100011010100110001010110001100011010111; end
            14'd408 : begin out <= 64'b0001111001100010000111011010100100100111111001111010100001011100; end
            14'd409 : begin out <= 64'b0010100011000001001001101001100000101010111101001010101100101110; end
            14'd410 : begin out <= 64'b1010101010000111001010011101010100101011010001111010100000101110; end
            14'd411 : begin out <= 64'b1010101111111111101010111010010010100111000101011010100100110101; end
            14'd412 : begin out <= 64'b0010100101010000001001001011000110101000000001011010100011110101; end
            14'd413 : begin out <= 64'b0001100110011011101010001010000010101010011110100010101011000010; end
            14'd414 : begin out <= 64'b0010101101111011101010110001010100100101010001111010101111111011; end
            14'd415 : begin out <= 64'b1000010000010110101000011011000110011111001010001010100111001111; end
            14'd416 : begin out <= 64'b1010000111011110101010010110100110101000100010110010010001010101; end
            14'd417 : begin out <= 64'b1010000111001001001001010000001000011010010111000010101111010100; end
            14'd418 : begin out <= 64'b1010101101000100000110110101000100101001101101111001111010101001; end
            14'd419 : begin out <= 64'b1010000101110110001001111010011110101011011010000010011001001110; end
            14'd420 : begin out <= 64'b1010010111000001001001011101000110101010010010101010100110101111; end
            14'd421 : begin out <= 64'b0001100101101000001010111000101010011001010100000010101010110010; end
            14'd422 : begin out <= 64'b1010101010000111001001111111100110100000001011001010010110011011; end
            14'd423 : begin out <= 64'b1010011110010110001010010011101000100100010100010001011111010111; end
            14'd424 : begin out <= 64'b1010011011000100001010100100111010100100011001100010101000011100; end
            14'd425 : begin out <= 64'b1010101000010110100111011011100110100001100100001010100001010101; end
            14'd426 : begin out <= 64'b1010101111110011001010110110110100101001100011101010101100110101; end
            14'd427 : begin out <= 64'b0001111011110101001010101101110000101000001110110010101111000011; end
            14'd428 : begin out <= 64'b1010100010111011001010000001111110101000101010101010100101100010; end
            14'd429 : begin out <= 64'b0010000110100100101010110101100010101000111001100010010010011000; end
            14'd430 : begin out <= 64'b0010100010000010101010000011110000101011111001101010101101011011; end
            14'd431 : begin out <= 64'b0010101110001000101010100010110110101001101110010010001001001101; end
            14'd432 : begin out <= 64'b1010101011111000100101111000001010101000101101000010100110011010; end
            14'd433 : begin out <= 64'b1010101000011011001000000010100000011101000110111010100101011011; end
            14'd434 : begin out <= 64'b0010100011101001001000110000101010101000011100001010101010111110; end
            14'd435 : begin out <= 64'b1001111110110110101001100111011110101000001101110010100101010011; end
            14'd436 : begin out <= 64'b1010100011011000001010110111001000100011101110110010000101111111; end
            14'd437 : begin out <= 64'b0010101100110001101010110110010010010111110001010010100111110101; end
            14'd438 : begin out <= 64'b1010011010010010001000001001000110101000000010111001101010100111; end
            14'd439 : begin out <= 64'b0010100000010000101001110011110110101001111111101010101011111101; end
            14'd440 : begin out <= 64'b0010000001011111101010110101011000101100000000101010100001000010; end
            14'd441 : begin out <= 64'b0010101000101110101001010110101010100111110101101010011011111000; end
            14'd442 : begin out <= 64'b1010100101111100001010001101111010100100010111010010101110000000; end
            14'd443 : begin out <= 64'b1010010100001111001010000100000000101000111001111001011110100101; end
            14'd444 : begin out <= 64'b1010101011101110100111100001001000100010110011110010000000100010; end
            14'd445 : begin out <= 64'b1010010100010010001010011100001100101010011010011010100101100101; end
            14'd446 : begin out <= 64'b0010010101111001101010001110000100101000001011101010000111010001; end
            14'd447 : begin out <= 64'b0001110001111110001010000110110100101001100101000010001111101000; end
            14'd448 : begin out <= 64'b1010101100001111100011100100011110100011101001110010010100100110; end
            14'd449 : begin out <= 64'b1001101111111001101010010111110100101010111100010010000101011011; end
            14'd450 : begin out <= 64'b0010010100011101101010101100000100101001110000000001111100100100; end
            14'd451 : begin out <= 64'b1010100011001010001010110001001100101010100010101010001001011100; end
            14'd452 : begin out <= 64'b0010001011100001001010110010000100101000100000011010100101010110; end
            14'd453 : begin out <= 64'b0010011101010001101010110001001010100111010000110010100001110101; end
            14'd454 : begin out <= 64'b1010100101101101100111011100000110011110111101011010010101101000; end
            14'd455 : begin out <= 64'b1001001010111110101010100010000000101001011001011010000111010111; end
            14'd456 : begin out <= 64'b0010001111111111101001011010101010101000010101110010100010011110; end
            14'd457 : begin out <= 64'b0010101010101101101010101110110110100100011010010010000110111110; end
            14'd458 : begin out <= 64'b1010101001000111001010111101101100101001100100011010101000000001; end
            14'd459 : begin out <= 64'b1010011111011001101010011110100010100110010100111010101100110110; end
            14'd460 : begin out <= 64'b1010011111100001100100010100001100100101001001000010011100011110; end
            14'd461 : begin out <= 64'b0010100111011010101010100100110100101001100111111001101010001100; end
            14'd462 : begin out <= 64'b1010001000011001100110011111010110101000111101111010100001001011; end
            14'd463 : begin out <= 64'b1010000011101101001010000101000000101011000111110010101101111001; end
            14'd464 : begin out <= 64'b1010010010010111001001111000001010100101010111110010000011110101; end
            14'd465 : begin out <= 64'b1001111101000010001001100010111000011011100101101010010010010000; end
            14'd466 : begin out <= 64'b0010001010110010001001101110010110010110100010110010101000001011; end
            14'd467 : begin out <= 64'b1010100111001011101010000010111000100111011101100010101010100100; end
            14'd468 : begin out <= 64'b1010100100101000101001000001001000101000000111100010100011100001; end
            14'd469 : begin out <= 64'b0010011011110101101001100101011010101010000011001010101110001111; end
            14'd470 : begin out <= 64'b0010010100001100101010011111010100010000001100100010101110111001; end
            14'd471 : begin out <= 64'b1010010011101100101010001100001000101010000100100010001111001110; end
            14'd472 : begin out <= 64'b0010100011110000101010011010100110011111100010101010101001100111; end
            14'd473 : begin out <= 64'b1010010001111110000101100111101010011010010000000010100000100100; end
            14'd474 : begin out <= 64'b0010011111011010101010001000010110101000000011100010101000101111; end
            14'd475 : begin out <= 64'b0010010110001001101001010011000000100011110111001010011100110000; end
            14'd476 : begin out <= 64'b0001111000010000100111111011001010101010000111101010100110101001; end
            14'd477 : begin out <= 64'b0010010101000100101010110001100100101000101101110001110101100100; end
            14'd478 : begin out <= 64'b0010101100110000001000101000100100101001110100101010010100011000; end
            14'd479 : begin out <= 64'b1010100100111011001001100100000110101000001100111010100001110100; end
            14'd480 : begin out <= 64'b0010010000011010101011000010001000101000001001000010010100000001; end
            14'd481 : begin out <= 64'b0010100110011100001010110111010000100100100001110010001000111000; end
            14'd482 : begin out <= 64'b1010001001010001101010111101010000101000101100111001111010010010; end
            14'd483 : begin out <= 64'b0010110000000010000011000010010000101001100110101010100000001001; end
            14'd484 : begin out <= 64'b0010011110000100101011000011001000100111010000010010101011100110; end
            14'd485 : begin out <= 64'b1010000001001011100110000010001100101010100001111010101111000010; end
            14'd486 : begin out <= 64'b1010100111010101001001001001010100101011101100011001110100001110; end
            14'd487 : begin out <= 64'b1010101000110101000111011110001000101000001111011010011010010000; end
            14'd488 : begin out <= 64'b0010100111110100001001001110100110101000001000011010011011010000; end
            14'd489 : begin out <= 64'b1010011001000010101001110111001010101001100010000010100010011100; end
            14'd490 : begin out <= 64'b0010010011011001101000011011111110101010001000001010101110000010; end
            14'd491 : begin out <= 64'b1010001100001100101010110100010100101001111111100010000110010000; end
            14'd492 : begin out <= 64'b0010011111111000101001001001110100100101000101011010100011111111; end
            14'd493 : begin out <= 64'b1010101010000011101010000000000100101010100001011010101000011100; end
            14'd494 : begin out <= 64'b0010010000011110001001110000001100101001000001000010101001110011; end
            14'd495 : begin out <= 64'b1010100011010000101010100010100110101010001111110010100011100111; end
            14'd496 : begin out <= 64'b1010100111100010101000101100001010100100010110100010100111000111; end
            14'd497 : begin out <= 64'b0010001101010101001010010111011000100010111001111010101101001010; end
            14'd498 : begin out <= 64'b1010100100100000101001011000011000101000100011010010011001000000; end
            14'd499 : begin out <= 64'b1010101000000001001001010010110010101001100000000010101011001010; end
            14'd500 : begin out <= 64'b1010100111111000001010000100100010101000000001001010010000010010; end
            14'd501 : begin out <= 64'b0010010100101110001010010110100100101000011010110010001000001101; end
            14'd502 : begin out <= 64'b1010100111110110100111101110100110101001111010011010101010101010; end
            14'd503 : begin out <= 64'b0001110110110001101010101011000100101001011001001010010111010001; end
            14'd504 : begin out <= 64'b0010000000011010101010001111110000101000000111111010000001010100; end
            14'd505 : begin out <= 64'b1010010001000100001010110110000000100100111111011010010110011000; end
            14'd506 : begin out <= 64'b1001110110100010101010100111101110101010101011010010001010111111; end
            14'd507 : begin out <= 64'b1001110100100101001001000001010100101100000010011010101111010001; end
            14'd508 : begin out <= 64'b0010101011011110001001010100111110100100010000110010011110101011; end
            14'd509 : begin out <= 64'b0010001010000110101010011010010000101010011111110010001010101101; end
            14'd510 : begin out <= 64'b0010100101111111101000101110010000101011101010000010100000100111; end
            14'd511 : begin out <= 64'b1010001011000010001010110011101000100100101100000001110101100000; end
            14'd512 : begin out <= 64'b1001101101000000100111001000010010100011100100010010001111000010; end
            14'd513 : begin out <= 64'b1010000010001010101000101110100100101001111111001010001110011111; end
            14'd514 : begin out <= 64'b1010100011000010101010110001010110101011011100000010010010010010; end
            14'd515 : begin out <= 64'b1010101100101111001010100000111010100100001000010010100001100001; end
            14'd516 : begin out <= 64'b0010100110110011001010101010011000011111010011100001000101001111; end
            14'd517 : begin out <= 64'b1010010000011101000111010011000110101011101101101010010110011100; end
            14'd518 : begin out <= 64'b0010100010110100101010001111001110010100101110011010100110100010; end
            14'd519 : begin out <= 64'b1010010001101011001010100111001100100110100110111010011001110000; end
            14'd520 : begin out <= 64'b0010001001001000001000101001101000100110101111111010101001111001; end
            14'd521 : begin out <= 64'b1010010111100000101010000100100100010110000101001010101111011000; end
            14'd522 : begin out <= 64'b1010101000101111000111110001100110101000001000100010011111011111; end
            14'd523 : begin out <= 64'b1010101101111010101000101101011100101010010000011001110110001010; end
            14'd524 : begin out <= 64'b0010100001110010001001101101101000100010001011100010101101001010; end
            14'd525 : begin out <= 64'b0010000010110111100111111000100100100100111100011001101011011100; end
            14'd526 : begin out <= 64'b1010100100010101100111000101111100100110110110010010010111110000; end
            14'd527 : begin out <= 64'b0001110110001001001010100010001000101001101110100010100011100101; end
            14'd528 : begin out <= 64'b0010101110010001001000000000110000101001010011011010011001100111; end
            14'd529 : begin out <= 64'b1010010011000100001001100101110110101010101111110010100101111111; end
            14'd530 : begin out <= 64'b1010100011100111101010011100010100100100100001001001011100011101; end
            14'd531 : begin out <= 64'b1001010101000010001010101111011000101011110000010010011111101111; end
            14'd532 : begin out <= 64'b0001101000000101101001010001100000101001010100000010100000000111; end
            14'd533 : begin out <= 64'b0001101100010111001010000010010010101000111100110010101001000011; end
            14'd534 : begin out <= 64'b0010000001010011001010011100100000100110011110110010101111001001; end
            14'd535 : begin out <= 64'b0010100100011110101010001000101000100010011000011010101010011001; end
            14'd536 : begin out <= 64'b1010010110110011101010101110111110101001011010010010101111111101; end
            14'd537 : begin out <= 64'b0010101011100101101010001111001000100101011010001010100011000101; end
            14'd538 : begin out <= 64'b0010101000101111001010100000000010100110101010100010010101011010; end
            14'd539 : begin out <= 64'b1010101011010001101010000001010100101000000010100010101110111000; end
            14'd540 : begin out <= 64'b0010000111100100101010101110110010011101011000100010100011001101; end
            14'd541 : begin out <= 64'b0010010111110010001001101001110110101011000011101010001010000010; end
            14'd542 : begin out <= 64'b1010100011001011001000001111111100101011110110001001110111100100; end
            14'd543 : begin out <= 64'b1010100111100011101001000110110100100101000101011010100100010010; end
            14'd544 : begin out <= 64'b0010001011001000001010110111110100101011011000111010011110100100; end
            14'd545 : begin out <= 64'b1010101001000111001000001101011110100111101011101010101000011001; end
            14'd546 : begin out <= 64'b0010101000001011101010101101010000100110101001100010101101001100; end
            14'd547 : begin out <= 64'b0010101001001101100111100111010100101011000110011010100010000000; end
            14'd548 : begin out <= 64'b0010010110010111001010100101011100100110010110110001110011010111; end
            14'd549 : begin out <= 64'b1010000010001001001010000001011100101001101000101010101101100110; end
            14'd550 : begin out <= 64'b1001000111100010101001111010101100100101001110001010101011110100; end
            14'd551 : begin out <= 64'b1010010111100011101001101010101000100011110100101001110110010011; end
            14'd552 : begin out <= 64'b0010100011110010001000101001010100100110110101110010100110011001; end
            14'd553 : begin out <= 64'b1010100101000000001010100111110010100110110100110001111100011101; end
            14'd554 : begin out <= 64'b0010001100000111001010010111011000100011110001000010000111111100; end
            14'd555 : begin out <= 64'b0001110010101011100110110011001010101001111010001010101111010110; end
            14'd556 : begin out <= 64'b1010100011010001101000101101000110101000101101010010010101100010; end
            14'd557 : begin out <= 64'b0010110000000001001000000000000010011110100101000001110110010110; end
            14'd558 : begin out <= 64'b1010011101010011101010101001010000101001110001101010010100010101; end
            14'd559 : begin out <= 64'b0010100011011110101001010111101010101011000010000010100011000111; end
            14'd560 : begin out <= 64'b0010000101010011001010110111110100100100010001011010100111110110; end
            14'd561 : begin out <= 64'b0010010000100001001010100000000110100010100000001010100101111000; end
            14'd562 : begin out <= 64'b0010011110110000100111000101001010100101000101001010000001111010; end
            14'd563 : begin out <= 64'b1010011100110011101010111001110000100110101110001010101010010011; end
            14'd564 : begin out <= 64'b1010101101001000001010101101101110101001101000100010101111100010; end
            14'd565 : begin out <= 64'b1010001100000010001001011110011110101001001001110010011100011001; end
            14'd566 : begin out <= 64'b0010100111000101001010010111011010101000010110111010101001101001; end
            14'd567 : begin out <= 64'b0010001100110110001010110110011110100110111111101010100110011111; end
            14'd568 : begin out <= 64'b0010101001001000001001011000010110100010011111101010100001000100; end
            14'd569 : begin out <= 64'b0010011001100001101001110111000010100101111000101010100111000001; end
            14'd570 : begin out <= 64'b1010101110100100001010111101001100011100111111001010011001001101; end
            14'd571 : begin out <= 64'b1010101011101001000101010010010100100111000111101001110100001100; end
            14'd572 : begin out <= 64'b1010011100010101101010001101001010100000100101000010100011101111; end
            14'd573 : begin out <= 64'b1010100010000010101010110000110010100111000111010001110010001000; end
            14'd574 : begin out <= 64'b1010100001001110001001101000011100100001001000101010000101011110; end
            14'd575 : begin out <= 64'b0000110000010111000111011001011010100111010000100010101001101110; end
            14'd576 : begin out <= 64'b0010011111000000101010001000011000100000000110001001001100100101; end
            14'd577 : begin out <= 64'b0010010001011110101010001011101100101001011100100001101100101000; end
            14'd578 : begin out <= 64'b1010000000011011101010000001001000100011010111111010101111110100; end
            14'd579 : begin out <= 64'b1001111111101110101010101101101100100001100001110010100111010101; end
            14'd580 : begin out <= 64'b0010101111011001100110101101100000101000111100111010100000111011; end
            14'd581 : begin out <= 64'b0010011101111100101001001100000010100111011001010010010001111010; end
            14'd582 : begin out <= 64'b1010010000001001000111010001111110101001011001110010011110011101; end
            14'd583 : begin out <= 64'b1010001011001000101000011101110110100110010010010001011000000110; end
            14'd584 : begin out <= 64'b1010101010000010001001001100111000101000001001000010100100011111; end
            14'd585 : begin out <= 64'b0010011111100100101001110001001010101010111011000010101100101000; end
            14'd586 : begin out <= 64'b1010101000100000001001110010110100101000110001011001011101000110; end
            14'd587 : begin out <= 64'b1010100101101000101010101100100000100001100101001010101111100101; end
            14'd588 : begin out <= 64'b0010100110000111101010101100001000011101101110000010001001101011; end
            14'd589 : begin out <= 64'b1010011100011100101001100110110010100011000000010010001010000011; end
            14'd590 : begin out <= 64'b0010011010000111101010011101010000100110001001111010000101110101; end
            14'd591 : begin out <= 64'b1010000011111010001010110110010110101010001110110010101101010110; end
            14'd592 : begin out <= 64'b0010100010000001001001001011011100101011110011000010101110101001; end
            14'd593 : begin out <= 64'b0010010111001001001001010101110000100110011011011010000101101010; end
            14'd594 : begin out <= 64'b1001011101111100001010110010000100011101011010101010100001010011; end
            14'd595 : begin out <= 64'b1010100100111010101001010111001000100001010110101010011001001110; end
            14'd596 : begin out <= 64'b0010001000101011101001010111001110100100010101100010100011110111; end
            14'd597 : begin out <= 64'b0010001010010000001010001111110010100000111110100010011010001000; end
            14'd598 : begin out <= 64'b1010011001000101101010110110100100011100110011010010010110000011; end
            14'd599 : begin out <= 64'b0010100110110110101010110000011110101001101101000010010111011111; end
            14'd600 : begin out <= 64'b0001111010000101101001001110010000101001110001110010100101110101; end
            14'd601 : begin out <= 64'b0010001111101101101010100111101010100010101101111001101010000001; end
            14'd602 : begin out <= 64'b0010100110011000100111001010110000101010110110110010100001100010; end
            14'd603 : begin out <= 64'b1010011100001010001000011110001100011010101011000001111101001000; end
            14'd604 : begin out <= 64'b0010011001001100101001011011111000011110111100100010100010011100; end
            14'd605 : begin out <= 64'b0010100110101110101000111010011010101001010100010010100001100001; end
            14'd606 : begin out <= 64'b1010100000010101100011111001111100010010010100000010101111001110; end
            14'd607 : begin out <= 64'b0010011111111000101010001101001110011101100101110010100011100110; end
            14'd608 : begin out <= 64'b0010010101010010000110001011100000100101101001100010100011110100; end
            14'd609 : begin out <= 64'b1010100110110101101000011110101000100100101011111010101100010110; end
            14'd610 : begin out <= 64'b1010001111010010101010010111010100100111010010111010100100110000; end
            14'd611 : begin out <= 64'b1010100111100000001010111011101110101011111101100010000111100110; end
            14'd612 : begin out <= 64'b1010001111110101001010011010000000011110011011011001100100111000; end
            14'd613 : begin out <= 64'b0010000110000111101010011011010110100010011011110010101011010101; end
            14'd614 : begin out <= 64'b0001101101011011100110000001011100101010011001001010010010101011; end
            14'd615 : begin out <= 64'b1010010101000001001010000110010010101010111011010010010000110000; end
            14'd616 : begin out <= 64'b0010010101100010101010101010011010101001011001100010100000110100; end
            14'd617 : begin out <= 64'b0010000101101010101001010110011000101011100101101001110111101011; end
            14'd618 : begin out <= 64'b1010101010011010001000100101110010101001010111101010010100000101; end
            14'd619 : begin out <= 64'b0010001101000010001010100111100110101010001100111010100101011011; end
            14'd620 : begin out <= 64'b0010101001110000101001010100010100100110110111110001111111010000; end
            14'd621 : begin out <= 64'b1010001010101011001010000100000000101010101001101010101011000111; end
            14'd622 : begin out <= 64'b1010100010101101101010111100011000101001111101011010100100111001; end
            14'd623 : begin out <= 64'b1010010010001111001010010010001010101001110111101010100011100011; end
            14'd624 : begin out <= 64'b1010100000001100101001010100011000100101011010000010010000110001; end
            14'd625 : begin out <= 64'b0010001101011111100101111110001000100110101110101000110111011110; end
            14'd626 : begin out <= 64'b1010101110000010101010001011010110101000100010101010000011000001; end
            14'd627 : begin out <= 64'b1010101100101100001000111100001000100001111010001010100110010001; end
            14'd628 : begin out <= 64'b0010010000011001101010110110110110101001100001101010100110111010; end
            14'd629 : begin out <= 64'b0010011111110111101010111100000110101011010100010010101101110011; end
            14'd630 : begin out <= 64'b1001010001110000101001110100101000101010011000011010011001011110; end
            14'd631 : begin out <= 64'b1010100000101100001000011001010110101011100101110010100001101110; end
            14'd632 : begin out <= 64'b1010101011101010000101011111001100101010110101000010000000110000; end
            14'd633 : begin out <= 64'b1010100111110101001010011101010010100001100111010010011010011001; end
            14'd634 : begin out <= 64'b0010101111100111001001100010001000101010010000010010010001011110; end
            14'd635 : begin out <= 64'b0010101101101011101010010011100100001110010010011010010100111010; end
            14'd636 : begin out <= 64'b0010101110100001101001000000101110100001010001010001011101100011; end
            14'd637 : begin out <= 64'b0010011111111010100111101110000100100111100011100001110001100000; end
            14'd638 : begin out <= 64'b0010100001010101001010001011011100101000101110001010101100000000; end
            14'd639 : begin out <= 64'b1010011001000111001010000000101110101001111110001010010101010000; end
            14'd640 : begin out <= 64'b0010011101000110101010100111100010100110010101000010100110100000; end
            14'd641 : begin out <= 64'b1010100111100100101010100111101000100110100111101010100010111001; end
            14'd642 : begin out <= 64'b0010000000011101101001111000000100011110001110010010011011000011; end
            14'd643 : begin out <= 64'b1010101110011001101010010000010110010001011110111010010100100111; end
            14'd644 : begin out <= 64'b0010011111111111101010010011010110100110010000001010100101000111; end
            14'd645 : begin out <= 64'b1010101010110110100111110010011010101010001000011010010011010101; end
            14'd646 : begin out <= 64'b0010101011110100001010011110001110011101001011000010100001000100; end
            14'd647 : begin out <= 64'b1010100001111101101000000010011110101011001001110010100101010001; end
            14'd648 : begin out <= 64'b0010010101011110101010101111111100101001001011001010010111111010; end
            14'd649 : begin out <= 64'b0001101001110100001001101010011010100101000100000010001101100100; end
            14'd650 : begin out <= 64'b0010001000011000100111011010101100101000000100111010101101011111; end
            14'd651 : begin out <= 64'b1010010010100111101010100100110000100100011010001010101001010011; end
            14'd652 : begin out <= 64'b0001111001110000100111010000100110010100101101110010011101110111; end
            14'd653 : begin out <= 64'b0010100011101001001010100010110100101001100000000010101110000101; end
            14'd654 : begin out <= 64'b0001110111110010001000000111101110100011000001111010000110001111; end
            14'd655 : begin out <= 64'b0010010011011011000111011110110110100110101100000010000101001111; end
            14'd656 : begin out <= 64'b1010100110111010000011110011111110101011010001000010100100010011; end
            14'd657 : begin out <= 64'b1010101100000001001001100110001000100011111110001010100000101000; end
            14'd658 : begin out <= 64'b0010100010010011101010010010110110101010111111011001101111101100; end
            14'd659 : begin out <= 64'b0010011010010000001010000100110000100101011001100010000000101001; end
            14'd660 : begin out <= 64'b0010001111100101001001000110001100101010101100100010011001110110; end
            14'd661 : begin out <= 64'b0010101011110001101000100010111110101010001101111001011011110110; end
            14'd662 : begin out <= 64'b0010011011101110101010001011001010011111001011010010101010000010; end
            14'd663 : begin out <= 64'b0001111101111000101001100100000110101000111001110010101011010101; end
            14'd664 : begin out <= 64'b1001111011010000100111010000001110100100011011101010101001000011; end
            14'd665 : begin out <= 64'b0010101101010010101000100111011110101000000010111010101010101101; end
            14'd666 : begin out <= 64'b0010100011001011001010100001101000101000010101100010010100101101; end
            14'd667 : begin out <= 64'b1010100110111000101001101010010100101000000001010010011001101001; end
            14'd668 : begin out <= 64'b1010101110100011101010010010111100100101101011010010011001000001; end
            14'd669 : begin out <= 64'b0010101001111111001001110101011100101000111100000010000110100011; end
            14'd670 : begin out <= 64'b0010011111001001001000101000001100100100000000011010101100001011; end
            14'd671 : begin out <= 64'b0010100110011000001010101001101100100111110111010010011111000011; end
            14'd672 : begin out <= 64'b1010100100000100001010110010000100101010011011001010000101111010; end
            14'd673 : begin out <= 64'b0001100110000011001010111010010010101001111001110001001001110000; end
            14'd674 : begin out <= 64'b1001010000111100001010111100011000101001010001001001110110100101; end
            14'd675 : begin out <= 64'b1001011100111101101001011110111010011101000000011010110000100101; end
            14'd676 : begin out <= 64'b1010000110100000101010011010100100101011100001110001101000100010; end
            14'd677 : begin out <= 64'b0010101101111111101001110111000010100000101110111010001010001010; end
            14'd678 : begin out <= 64'b1010100011100011001010111111000100101000011010110010100100110100; end
            14'd679 : begin out <= 64'b0010101000100010101010110110000000101001001110111010100101111110; end
            14'd680 : begin out <= 64'b0010101011011101001001101010011010101000101001101010101101011001; end
            14'd681 : begin out <= 64'b0010001000101001001010011010110100100100010011100010011100001111; end
            14'd682 : begin out <= 64'b0010010100110100001010100101101000101011000011110010101000110011; end
            14'd683 : begin out <= 64'b0010011111100000101010001000101100100010000000101001000100111011; end
            14'd684 : begin out <= 64'b1010101011111001101010001010110100101001010100101010100000100000; end
            14'd685 : begin out <= 64'b0010000101101100001000101110101110100010110001010010001000000011; end
            14'd686 : begin out <= 64'b1010000111000011001001100111101010101010010101101010100010001001; end
            14'd687 : begin out <= 64'b0010011111001100101000101111100100100100000010001010011100110000; end
            14'd688 : begin out <= 64'b1010100011110010101010110011011100101000011010001010001010101101; end
            14'd689 : begin out <= 64'b0010001100111110101010101011011010101001001011000010101001100011; end
            14'd690 : begin out <= 64'b0010000010101010101000011110011010011001110010000010100010011100; end
            14'd691 : begin out <= 64'b0010101110100110001010011011000100101000111001011010101000000010; end
            14'd692 : begin out <= 64'b1010010101011000101001001101100000101010011011010010011010001101; end
            14'd693 : begin out <= 64'b1001011100101001001001100111100100101011010001111010001101011000; end
            14'd694 : begin out <= 64'b0010100000001100001010100010111110101000011100010010010001111110; end
            14'd695 : begin out <= 64'b1010000010011110101001010001010000101011000101000010000101000000; end
            14'd696 : begin out <= 64'b1010101001010000101010111000010100100100101100000010100101001111; end
            14'd697 : begin out <= 64'b1010011010001110001010000001010110101001010011111010011010111110; end
            14'd698 : begin out <= 64'b0010001111110000101010000010100010100100010001010010010011111111; end
            14'd699 : begin out <= 64'b0010101001101010000111010100010010101010000110011010101101011011; end
            14'd700 : begin out <= 64'b1010011111010001100111111111111100100100000100111010100000110101; end
            14'd701 : begin out <= 64'b0010101011110001101010000100011110100100101100111010101100110000; end
            14'd702 : begin out <= 64'b1010010010100110101001010011011000101001000111001010100110110010; end
            14'd703 : begin out <= 64'b1010101001110101101001000001101000011000101111000010000011111100; end
            14'd704 : begin out <= 64'b0010101011010000001010000101100110101000111110101010100001110010; end
            14'd705 : begin out <= 64'b1010101111000000001001010110010010101000000110111010000111101111; end
            14'd706 : begin out <= 64'b0010101110001010101001100110111000100110010001001010011000011011; end
            14'd707 : begin out <= 64'b1010100101111111001001110101001000101010100001011010000111101011; end
            14'd708 : begin out <= 64'b1010100101000101001010001000010100011100000010111010011010110000; end
            14'd709 : begin out <= 64'b0010100101000001001010000101001000011011100001001001010100101011; end
            14'd710 : begin out <= 64'b0001100110111000000110110101010010101001110111110010100010000000; end
            14'd711 : begin out <= 64'b1010011000101011001010101100110010101011011111001010011000010110; end
            14'd712 : begin out <= 64'b0010010100110101101010010011001000101001101010101010010100111111; end
            14'd713 : begin out <= 64'b1010101011000101001010110100101100011110010101110010010100001101; end
            14'd714 : begin out <= 64'b0010100111111101101010000110100100101011011010001010101010001101; end
            14'd715 : begin out <= 64'b0010101101000101101010010110011100100111000110010010000001011001; end
            14'd716 : begin out <= 64'b1010010111100111000111110111000100101001010010100010101010100011; end
            14'd717 : begin out <= 64'b1001001000001110001010000101001010100110010011111010100011111100; end
            14'd718 : begin out <= 64'b1010011101111000101010110010100110100101011101101001100101100011; end
            14'd719 : begin out <= 64'b1010101011111111101010011100111100101001101111011010101111011010; end
            14'd720 : begin out <= 64'b1010100101000000001010011101111010101011111011111010100010011111; end
            14'd721 : begin out <= 64'b0001111100011010101010111001011100100110011010110010000001111100; end
            14'd722 : begin out <= 64'b0010011111011101001010111111110110011010001101101010101010000101; end
            14'd723 : begin out <= 64'b0000110001100010001000010001010000101011011011100010000101111010; end
            14'd724 : begin out <= 64'b0010100011110000001001000110111000100101100000111010010110011111; end
            14'd725 : begin out <= 64'b0010101001011111101001101001110010100111000010100010101101000010; end
            14'd726 : begin out <= 64'b0010000110000001001010110101100100101001001100110010101010011101; end
            14'd727 : begin out <= 64'b0010011111100110001010000000101100101000110110110010100100001010; end
            14'd728 : begin out <= 64'b0010100101010010001001001110010010100101011101101010000111000011; end
            14'd729 : begin out <= 64'b1010101001010110101010000111110000100110100111010010011000111100; end
            14'd730 : begin out <= 64'b1010101111011110101001001011111100101000010000100010101101110111; end
            14'd731 : begin out <= 64'b1010100011000111101000110011110100101011000110111010011001010110; end
            14'd732 : begin out <= 64'b1010000100101100001010100011100110100100010010011010011100001011; end
            14'd733 : begin out <= 64'b0010011011111011000101101100111000101010100110000001111110100111; end
            14'd734 : begin out <= 64'b1010011111010011001010010001001010101011101111001010101011100000; end
            14'd735 : begin out <= 64'b1010000000111000100111011101111000101000111100111010100010111101; end
            14'd736 : begin out <= 64'b1010100010000100001010101000001100101001100000000010011001011000; end
            14'd737 : begin out <= 64'b0001100111010010101010100100000100101010011000001010001010101001; end
            14'd738 : begin out <= 64'b1010001010101100101010110100110000100111010111110001110000100100; end
            14'd739 : begin out <= 64'b1010101100111000001010100011100110101010100110001010010101011011; end
            14'd740 : begin out <= 64'b0010101000101110100111010100000110101001011101110010101111100110; end
            14'd741 : begin out <= 64'b0010011110111011001000101100011100001110010100101010001100001100; end
            14'd742 : begin out <= 64'b0010100010000000001001011011111100101011111011110010001001011101; end
            14'd743 : begin out <= 64'b0010101101111010001010000101011010011100101010101010100111110101; end
            14'd744 : begin out <= 64'b1001111101011001101000110011011010100101011101110010011111111011; end
            14'd745 : begin out <= 64'b0010100110010111101010001001110100100101100000000001110110110011; end
            14'd746 : begin out <= 64'b1010101010011101001001111101010100100101011000010010001010111011; end
            14'd747 : begin out <= 64'b1010101100000101101000000011101000101001111100011010101010100100; end
            14'd748 : begin out <= 64'b1010010011101101001000100111000010100100111000110010011011001001; end
            14'd749 : begin out <= 64'b0010101000110000001010000100010110100111010011011010011101110101; end
            14'd750 : begin out <= 64'b1001101100010101100111110100000010101011001000000010101111101100; end
            14'd751 : begin out <= 64'b0010101010101100101001010011010000101010110001000001110110010001; end
            14'd752 : begin out <= 64'b1010011111110110001000011100100000101011010011100010100000010100; end
            14'd753 : begin out <= 64'b0010101101001100101010010011011010100001101100001010011110101000; end
            14'd754 : begin out <= 64'b1010010001010000101000011001000000101011010110010010001101101001; end
            14'd755 : begin out <= 64'b0010101001100101101001010001100100100110110011011010100000111110; end
            14'd756 : begin out <= 64'b0010100100100010001010100000010000100011011111011010001100001100; end
            14'd757 : begin out <= 64'b1010011000101110101001110111111000101001110011100010011110101000; end
            14'd758 : begin out <= 64'b1010101000000100101000000001110110101011011010101010101000010010; end
            14'd759 : begin out <= 64'b1010010111111001101001010110111100101011101001100010100111000010; end
            14'd760 : begin out <= 64'b0010010100001100101001000001010100011010111100101010001110101100; end
            14'd761 : begin out <= 64'b1010101001010100100110101001111110011110011110000010101011011110; end
            14'd762 : begin out <= 64'b1010101001111101001000001110110110101000110000100010100111101110; end
            14'd763 : begin out <= 64'b0010101000110000101010011011000010100101010001101010101111100000; end
            14'd764 : begin out <= 64'b1010011011100000101010111111000110011111011000111010101101111101; end
            14'd765 : begin out <= 64'b1010100000100000101010100000000010011110111111001010010110111001; end
            14'd766 : begin out <= 64'b0001010010101001001010011000100100101000101010011010101000000010; end
            14'd767 : begin out <= 64'b1001101101011110001010100000111100101010011010100010100110110110; end
            14'd768 : begin out <= 64'b0010101011111000001010100010000110100100111101110010001011000001; end
            14'd769 : begin out <= 64'b0010011111100111000110001001001100011001100011101010000001110011; end
            14'd770 : begin out <= 64'b1010100010101100101001001100100110101010100110101010001100011101; end
            14'd771 : begin out <= 64'b1010011001101100001010010010010000100000111101111010010000000010; end
            14'd772 : begin out <= 64'b0010101111101001001010000011001000100110011001110010010100110111; end
            14'd773 : begin out <= 64'b1010011011111000101000000110010110101011100001110010101001101001; end
            14'd774 : begin out <= 64'b1010011101011110001010111010111100011111111000110010101110110010; end
            14'd775 : begin out <= 64'b1010101111001101001000111110011110101011010000011010100100010010; end
            14'd776 : begin out <= 64'b0010100000011000001010100111111000101000111010011010100110100001; end
            14'd777 : begin out <= 64'b0010100001111101001000011011111110101010001010010010000000011110; end
            14'd778 : begin out <= 64'b0010011001001000101010000101001110101011010010011010100100010001; end
            14'd779 : begin out <= 64'b0010000011011001101010011001010110100110100100000010100110100011; end
            14'd780 : begin out <= 64'b0010011110000100101001100111000100100110100001011010100011111000; end
            14'd781 : begin out <= 64'b1010010010100010000101010110011010011100111100011010001000110001; end
            14'd782 : begin out <= 64'b1010000001001111001010111001101000100000101111000010001001111011; end
            14'd783 : begin out <= 64'b1010101000110000001010101100010000101000100110011010101011110111; end
            14'd784 : begin out <= 64'b1010011110100000001010100101110000101010110111000010100001111011; end
            14'd785 : begin out <= 64'b1010101110011101101010001101111000100110111111001010101011101110; end
            14'd786 : begin out <= 64'b1010100011110010100111100001010000101000110000111001011011010000; end
            14'd787 : begin out <= 64'b0001011011111111101001001111101010100101000000100010011000100110; end
            14'd788 : begin out <= 64'b0010010011010100001010101011000010101000011101110010100110010001; end
            14'd789 : begin out <= 64'b1010000011111010001010100010111110101010100001010010101010001101; end
            14'd790 : begin out <= 64'b1010011001111101001001001011000110101000110101100010100010001110; end
            14'd791 : begin out <= 64'b1010101111001111001001100100101010101011011011111010001001111011; end
            14'd792 : begin out <= 64'b0010100000111011001010001001010000101010110000100010100101110111; end
            14'd793 : begin out <= 64'b1010011000101110001010000110100100101000101010010010000001100000; end
            14'd794 : begin out <= 64'b0010101000110011101000100100110000101011010101000010001111111000; end
            14'd795 : begin out <= 64'b0010100010011011101001001001010100101001110100001010100110101111; end
            14'd796 : begin out <= 64'b0010000100110010100111100101111110101001111001001010101001001100; end
            14'd797 : begin out <= 64'b0010101010000111101000101100101100101011000000010010100010001011; end
            14'd798 : begin out <= 64'b0001110101110000101000000000110100100010001011110000111100111100; end
            14'd799 : begin out <= 64'b0010101000000010001010101011101000100111100001000010100111110001; end
            14'd800 : begin out <= 64'b1010100011010000001001101110111100101010001101000010010011011111; end
            14'd801 : begin out <= 64'b1010010001011011001000001011001110101100000010100010101001011010; end
            14'd802 : begin out <= 64'b0010101000000000101001111110110110101010001011111010011011100011; end
            14'd803 : begin out <= 64'b0010000011100101101010011101100010100110110101100010100010111100; end
            14'd804 : begin out <= 64'b0010101000011111101001101010100110100101001000111010100100100010; end
            14'd805 : begin out <= 64'b1010100111100100101010010110111110011100110110111010010100101110; end
            14'd806 : begin out <= 64'b1010100110101000101010100111010100101010111011000010010111001001; end
            14'd807 : begin out <= 64'b1001010011111001101010011101110000100100100001111010101000011010; end
            14'd808 : begin out <= 64'b0010100110100000001001101001111000011110100101011010101101001000; end
            14'd809 : begin out <= 64'b0010011111100000001010110011101010101011001111110010100100001011; end
            14'd810 : begin out <= 64'b1001111000010110000111000011000110100110110101000010101000010101; end
            14'd811 : begin out <= 64'b0010001001010010001000010110010010011100011000011010011110100011; end
            14'd812 : begin out <= 64'b0001101101011010000110011110011110101001111110111010101011110001; end
            14'd813 : begin out <= 64'b1010010111110100001010110011100110100110010011101001111110011011; end
            14'd814 : begin out <= 64'b0010000010001110101001110000000110101010100010110010100101101001; end
            14'd815 : begin out <= 64'b0010101010011011100110101011010010100110110110101001011011001011; end
            14'd816 : begin out <= 64'b0010010111100110001010111001010110011110100001110010100101000111; end
            14'd817 : begin out <= 64'b0010101000100001001010010001010110101011000100000010010010011001; end
            14'd818 : begin out <= 64'b1010100010001100101010010001111110100111111001110010011101111010; end
            14'd819 : begin out <= 64'b0010001100001111001010000000100110100011000011111010010000011110; end
            14'd820 : begin out <= 64'b1010100110100111001000110011101010101000001000101010011100010000; end
            14'd821 : begin out <= 64'b1010100110100110001010101101001110100110101101011010101011001101; end
            14'd822 : begin out <= 64'b1010100011001111101001101000010000101010010111010010000100110101; end
            14'd823 : begin out <= 64'b0010101000011111001001111100101010101001011100110010100011101111; end
            14'd824 : begin out <= 64'b0010000100010001101001000101000100101011110101100010100011111101; end
            14'd825 : begin out <= 64'b1010101101110010001001010000011010100110001101011010100000110110; end
            14'd826 : begin out <= 64'b1010100001001001101001001000110110101001001011000010101001110001; end
            14'd827 : begin out <= 64'b1010101000011101001010001100111100101000101101110001101011001000; end
            14'd828 : begin out <= 64'b1010101000000111001010101011001010100110011000110010100101111011; end
            14'd829 : begin out <= 64'b0010101011111101101010011001011000011101100101010010001000011100; end
            14'd830 : begin out <= 64'b0010001100101111001010000110011000101010000100101010001111111100; end
            14'd831 : begin out <= 64'b0010100110000100000110011110111000101010001100111010000011101111; end
            14'd832 : begin out <= 64'b0010101010001010000101010110111100011110001100100010101010010111; end
            14'd833 : begin out <= 64'b1001111101000100001010110110100110101000110001010001110101110111; end
            14'd834 : begin out <= 64'b1010011110011001101000001111010010100101011010110010100111010110; end
            14'd835 : begin out <= 64'b1010010011100101001000000110000000011010010100110010101001111010; end
            14'd836 : begin out <= 64'b1010100010000010001010110011010100100000010101011010010100111110; end
            14'd837 : begin out <= 64'b0010001001111110100111101000001100101001111110111001100011100110; end
            14'd838 : begin out <= 64'b0001110011101010101010100101011100101010110110111010101101011010; end
            14'd839 : begin out <= 64'b0010100110000101001010011011000110101001100000001010001011101000; end
            14'd840 : begin out <= 64'b1010100100000011101001001000111100101001011000110010011001100100; end
            14'd841 : begin out <= 64'b1010100101001001001010100011010110100001100011000010101100101010; end
            14'd842 : begin out <= 64'b1010100001000000101001011101111010101010010100101010100010000001; end
            14'd843 : begin out <= 64'b1010100001101011001010111001100100101011110001111010100000111100; end
            14'd844 : begin out <= 64'b1010100000110100101001000100100000101001001101001010101000011110; end
            14'd845 : begin out <= 64'b0010100011010000001010110010111010101010111011001010100010111110; end
            14'd846 : begin out <= 64'b1010010111010011101010101111101100101001110000010010100011110100; end
            14'd847 : begin out <= 64'b0010001111010001001010001101001110101011100011010010101101010110; end
            14'd848 : begin out <= 64'b1010101011011111001010110111001000100101101010001010100001111110; end
            14'd849 : begin out <= 64'b0010010000100100101010000001001010101011001110100001110000000000; end
            14'd850 : begin out <= 64'b0001110101101101101010101000110100100100100000000010100110100011; end
            14'd851 : begin out <= 64'b0010010010110100001000001001101010100000000000110010100100011010; end
            14'd852 : begin out <= 64'b0010000100001111100110110011110110101011101101110010011110101010; end
            14'd853 : begin out <= 64'b1010101101000111101010011101010100100111100010111010010000110110; end
            14'd854 : begin out <= 64'b1010100011111100101001100101010100100011111011011010011110100101; end
            14'd855 : begin out <= 64'b0010001100010101001000010110000000101000011010011010011010101110; end
            14'd856 : begin out <= 64'b0010101111111011101010010111011000100001000001111010011100110111; end
            14'd857 : begin out <= 64'b0010011100000100101001111110010110100111110011101010101100001110; end
            14'd858 : begin out <= 64'b1010100111000000001000001110100010100101001001100010100111101110; end
            14'd859 : begin out <= 64'b1010000001101110001001000011100000101010001011010001111100001110; end
            14'd860 : begin out <= 64'b1010011111010000101010110001110000100110110110000010001110011111; end
            14'd861 : begin out <= 64'b0010000011000101101010011100001100100111101001100010100001011111; end
            14'd862 : begin out <= 64'b0010011100111101001010010001100000011101111110001010101001101010; end
            14'd863 : begin out <= 64'b1010100101001011101000010010100100101000001100111010100001010001; end
            14'd864 : begin out <= 64'b0010001111110001001010010100000100100010111111000010100010001100; end
            14'd865 : begin out <= 64'b0001100011010000001010011000011110011100101000000001110111111101; end
            14'd866 : begin out <= 64'b0010101000000010101010110100000010101010100110111010100001110010; end
            14'd867 : begin out <= 64'b1010101011010111001010101100101100100110001100101010001001101100; end
            14'd868 : begin out <= 64'b1010010001000110001010101101000000101000101110000010100011101010; end
            14'd869 : begin out <= 64'b0010101110110000101010001100110100101000001100100010100111001001; end
            14'd870 : begin out <= 64'b0010011010111000100101100111111100101001100110011010100000110000; end
            14'd871 : begin out <= 64'b1010101101011010001010110110011010100110110100010010100100011011; end
            14'd872 : begin out <= 64'b1010010011111000001000001110110010100100011011101010011110011110; end
            14'd873 : begin out <= 64'b0010001010100011001001111011011100100110000000111010101010111001; end
            14'd874 : begin out <= 64'b0010101101001101001010110100111110101010000000111010011111111100; end
            14'd875 : begin out <= 64'b1000110011010011101000101101111000101001101010001010100010010111; end
            14'd876 : begin out <= 64'b0010100011000100001000100100111010100110010011101010101110000000; end
            14'd877 : begin out <= 64'b0010010111100110000110100111001010101011100001011010101111101110; end
            14'd878 : begin out <= 64'b0010101011100000100100010101010110101000110010000010000101110111; end
            14'd879 : begin out <= 64'b0010010011110011101010100110010000011100111011011010101100110111; end
            14'd880 : begin out <= 64'b1010001010000101000001000011100000101001111111101010101111110001; end
            14'd881 : begin out <= 64'b1010011000010110101000111100111110100100011101111010010001000010; end
            14'd882 : begin out <= 64'b0010000111010010001010111110110010101000000011100010100100100001; end
            14'd883 : begin out <= 64'b0010101110101101101001111110100110100110001010000010101101000000; end
            14'd884 : begin out <= 64'b1010101111001110001001111111010010010001000001010010011110001111; end
            14'd885 : begin out <= 64'b0010010000101100101010111111001110101001001001101010101101110011; end
            14'd886 : begin out <= 64'b0010000010100111001010101100100000100000001010010010101001000111; end
            14'd887 : begin out <= 64'b0010100011111010101000010001001000101010001111100010011000100011; end
            14'd888 : begin out <= 64'b1010001010110111100110100101011000101000101101000010100100100010; end
            14'd889 : begin out <= 64'b0010101100100111101010010110101110101000101101010001110111010100; end
            14'd890 : begin out <= 64'b0010100001000110001001100001100110011001110001100010100000100000; end
            14'd891 : begin out <= 64'b0010100001101111001001011010101100101010001111110001111011111000; end
            14'd892 : begin out <= 64'b1010011011010101101000011100111110100001101101000001110010011100; end
            14'd893 : begin out <= 64'b0010100000110110001001011110001100101000001010110010100001100100; end
            14'd894 : begin out <= 64'b1010100011100010101010110101011000101011010010010010011000000100; end
            14'd895 : begin out <= 64'b1010010001011110101010001010101100101010010010011010100000110010; end
            14'd896 : begin out <= 64'b0010001011001110001000001001110100010111111000101010010010100000; end
            14'd897 : begin out <= 64'b1010100111000111101010011011010100011011000000000010101001110000; end
            14'd898 : begin out <= 64'b1010100010001010101000011001001100100110111000110010100010100000; end
            14'd899 : begin out <= 64'b1001110101010111101010100010000110011100010110100010100111010010; end
            14'd900 : begin out <= 64'b1010011111110001001010111011000110100100010001010010010000001100; end
            14'd901 : begin out <= 64'b1010010001100001001001110111001110100100011011010010101100001010; end
            14'd902 : begin out <= 64'b0010001110111011101010010111100010010100000100100010101001101010; end
            14'd903 : begin out <= 64'b1010011010001110101010110001100000101011000010111010001111100110; end
            14'd904 : begin out <= 64'b0001001100000001001000101010100000011111101010010010010111010000; end
            14'd905 : begin out <= 64'b1010101101111000001010000010010110100101011001110010100100001010; end
            14'd906 : begin out <= 64'b0010100010010000101010001101110010101011111110111010100010110010; end
            14'd907 : begin out <= 64'b1010011101000100001001101111101010010101001010001010011110000111; end
            14'd908 : begin out <= 64'b0010100000111110001010111011000100100101111001001010000010100000; end
            14'd909 : begin out <= 64'b1010000110101000001010011000011110100000101001010001111000001001; end
            14'd910 : begin out <= 64'b0010100001001110101010001010011010100001001000110010101100010000; end
            14'd911 : begin out <= 64'b1010101110011010101010110001101010100110100111000001110011101001; end
            14'd912 : begin out <= 64'b0010101111010001001001011111001010101000011010101010000011101011; end
            14'd913 : begin out <= 64'b0010011011001001101000011101100000101010011110110010100010101111; end
            14'd914 : begin out <= 64'b0010000000101010000111111111100010100001100101000010101001010000; end
            14'd915 : begin out <= 64'b1010011111111110001010011001000000100010110000010010100000101110; end
            14'd916 : begin out <= 64'b0010010000111010101010100111100100101010111101111010010111101110; end
            14'd917 : begin out <= 64'b1010101111110111001000101011100110100011100110101010010001111000; end
            14'd918 : begin out <= 64'b0010010000110110001010100111110110101011101101110010000110001010; end
            14'd919 : begin out <= 64'b1010100010011100101010110011111000011101010111100001110011010101; end
            14'd920 : begin out <= 64'b0010010111001111101001011101001110011101000010011010100011110111; end
            14'd921 : begin out <= 64'b0010010001011010000110111010011000100000011011100010100101111010; end
            14'd922 : begin out <= 64'b1010011010110111001010111010101010101011001000000010101010101110; end
            14'd923 : begin out <= 64'b0010100111010010001010010011111100100100111010100001110100100101; end
            14'd924 : begin out <= 64'b0010100100000010101000010000101000101001001101001010011000001001; end
            14'd925 : begin out <= 64'b1010100110111001101010010011010100100100111011111010101111110000; end
            14'd926 : begin out <= 64'b1010101001011010000110110110000100101010100001001010101010101001; end
            14'd927 : begin out <= 64'b0010011011000010100111001111100110101000011011110001111100010000; end
            14'd928 : begin out <= 64'b0010011010100011101010110000011000101010100101110010011011101111; end
            14'd929 : begin out <= 64'b1010010001101001101010101111001110100101110001100010101111001010; end
            14'd930 : begin out <= 64'b1010011100001111101010100010001000100111001101110010100001000110; end
            14'd931 : begin out <= 64'b1010100100110011101010101110101100011110101100000010010010011001; end
            14'd932 : begin out <= 64'b0001100110110010101010000101001000101011011001101010000010111101; end
            14'd933 : begin out <= 64'b1010101000111101101010111010010110100011000110110010100111101100; end
            14'd934 : begin out <= 64'b1010011111000100101001100101000000100101011111011001111101010100; end
            14'd935 : begin out <= 64'b0010100010110000001010100100110010100100101001111010101000011101; end
            14'd936 : begin out <= 64'b0010100110111001001001010100011110100100010111111010011001001101; end
            14'd937 : begin out <= 64'b1010101001001110001010110001110110101010101111100010011001001000; end
            14'd938 : begin out <= 64'b0010101111000110001010111011100010101010000010011010100100111110; end
            14'd939 : begin out <= 64'b0010010001001011001010000000000000101000101011000010010010010110; end
            14'd940 : begin out <= 64'b1010101000111110101001110011101100100100001000110010001001010000; end
            14'd941 : begin out <= 64'b0001100101001000001010101010111110100101100010001010101100100001; end
            14'd942 : begin out <= 64'b1010000110011100100111000111001000100001011101110010101010111111; end
            14'd943 : begin out <= 64'b0010101111011010001010100101110010101011000110001010100010101111; end
            14'd944 : begin out <= 64'b0010101100010000101010110010110100101011011110000010100011011100; end
            14'd945 : begin out <= 64'b1010101101001011001000001110111010101011101001111010011011100010; end
            14'd946 : begin out <= 64'b1001010001010011000111101101010000101010110111111010000100001000; end
            14'd947 : begin out <= 64'b1010101010111111101001011011011100101011101010111010001110000100; end
            14'd948 : begin out <= 64'b1010101000011110001010001010011010100101001011110010101100010010; end
            14'd949 : begin out <= 64'b0010001101101010100111010111011100100011001011110010000100100100; end
            14'd950 : begin out <= 64'b1010101111001100000100101100001100100100101110001010010000101110; end
            14'd951 : begin out <= 64'b1010101000001101001001101111010110100111101001010010100011011010; end
            14'd952 : begin out <= 64'b1010000111111010100101110011010010101011000001111010100010010001; end
            14'd953 : begin out <= 64'b0001110001100111101000111111000010100010100001100010100011110100; end
            14'd954 : begin out <= 64'b0010100011111101001001001111011010101010100011111010101111100001; end
            14'd955 : begin out <= 64'b0010101010001010001010110000100000100101100111010010010010101001; end
            14'd956 : begin out <= 64'b0010011101010101001010100010010010101001101101011010101101011000; end
            14'd957 : begin out <= 64'b1010001101110000001000010101001010101001011010010010101111010111; end
            14'd958 : begin out <= 64'b0010101010110011001010011011011110101010101110101001111111000101; end
            14'd959 : begin out <= 64'b0010010011100111101001100101001010101000000011011010100111001000; end
            14'd960 : begin out <= 64'b1010100001111010101010001110111110101001010110110001110011011011; end
            14'd961 : begin out <= 64'b1010000111111111101010000001100100101011110101000010010100011110; end
            14'd962 : begin out <= 64'b0001101100100100001010010111101100100001110010100010101101011111; end
            14'd963 : begin out <= 64'b0001100101101010101010111011000010100011001001101010101000011001; end
            14'd964 : begin out <= 64'b1010100111101000101010010001100100101011000000010001111000000110; end
            14'd965 : begin out <= 64'b0010100111000000100111011011100000101010101000010010000010111100; end
            14'd966 : begin out <= 64'b1001100101111111101010011111001010101011010000111010100011011110; end
            14'd967 : begin out <= 64'b0010010001110111101010101000011110100000111111100010001010011111; end
            14'd968 : begin out <= 64'b0010100001101110100101110101010100101001100000011010101000100011; end
            14'd969 : begin out <= 64'b0010010000101111001010000011000110101000011101100001111011010101; end
            14'd970 : begin out <= 64'b1010100100000110101000100100001000100111101010011010000101100001; end
            14'd971 : begin out <= 64'b1010001000011111000111110000001100100100010010101001110100010011; end
            14'd972 : begin out <= 64'b0010101110011101001010010100000100011000101111100010100111101000; end
            14'd973 : begin out <= 64'b0001111110110001101010011101000110101011011010010010101110001110; end
            14'd974 : begin out <= 64'b0001101110111111001001111010010010101011011011000010101101101100; end
            14'd975 : begin out <= 64'b1010010111011101101010010101011110101001011100110010010000011100; end
            14'd976 : begin out <= 64'b0010100011011000001010010110101010101011111000100010101100011001; end
            14'd977 : begin out <= 64'b1010101111111001001010001101100110100100111001111010101010000101; end
            14'd978 : begin out <= 64'b0010101001010000101001100101111010101000001011110010010111010110; end
            14'd979 : begin out <= 64'b0000111100011111000111100110111100101001000101111010101101001001; end
            14'd980 : begin out <= 64'b1010011100011111101001010110001010010110111101000010000100111111; end
            14'd981 : begin out <= 64'b0010001110000110000100010101110010100000001101010001100000111001; end
            14'd982 : begin out <= 64'b0001101011100001100111000001101110101011000001001010100111000010; end
            14'd983 : begin out <= 64'b1001100111111001001010011010111000101011010100000010100000011111; end
            14'd984 : begin out <= 64'b1010101111110011100101000101110110100111010100010010010110000001; end
            14'd985 : begin out <= 64'b0010001110000111101001100010100010100110001101101010101000100110; end
            14'd986 : begin out <= 64'b1001100000100011101000011100000110011111111101000001101110100011; end
            14'd987 : begin out <= 64'b0010101001111101001001011111011100100100100100011010000001000111; end
            14'd988 : begin out <= 64'b1010001111001010001001101100000010100111111100110010010010010101; end
            14'd989 : begin out <= 64'b0010100110000110101010010111001110100101000011010010011011000000; end
            14'd990 : begin out <= 64'b1010100000010000001000011110010000101010011011110010000100110001; end
            14'd991 : begin out <= 64'b0001100001111000001010101001011110100000100100011001011011111010; end
            14'd992 : begin out <= 64'b1001101101110101001010111101101100101000111101010010010000111111; end
            14'd993 : begin out <= 64'b1010011011110100101001100111011100101011100001101010010000010000; end
            14'd994 : begin out <= 64'b1010100000001101001010110110000100100110100011001010001100000110; end
            14'd995 : begin out <= 64'b0010100100011001101010001011101110100101101000101010101110101111; end
            14'd996 : begin out <= 64'b0010010101011101001000111101010100101010110111001010011111100110; end
            14'd997 : begin out <= 64'b1010000111111101101010110110000000100000010011010010101010011001; end
            14'd998 : begin out <= 64'b1010101011001010001001011001010100101000101110011010001101110001; end
            14'd999 : begin out <= 64'b1010001001000001101001011110110110101000010001100010011001111000; end
            14'd1000 : begin out <= 64'b0010011010110100000101010010110100010101110001110010010001111100; end
            14'd1001 : begin out <= 64'b0010011110010011101001101111010010001000001100100010011000001011; end
            14'd1002 : begin out <= 64'b1010101010001001001010011000011100100111111101010010101110011101; end
            14'd1003 : begin out <= 64'b1010011010101110101000111000010000100110001000001010101100000010; end
            14'd1004 : begin out <= 64'b1010101100110101000100100010001010101011110110010010101111100111; end
            14'd1005 : begin out <= 64'b1010100101001011101010111000101110101011110110000010100100010111; end
            14'd1006 : begin out <= 64'b0010100110001000001001101100010000101001010011010010101100000110; end
            14'd1007 : begin out <= 64'b0010101000100111101010101110000100101011100111100010011000010000; end
            14'd1008 : begin out <= 64'b0010101110110111101001011010101100101000000110111010101101111110; end
            14'd1009 : begin out <= 64'b1001110001101010101010111000101100100001000001101010011010011010; end
            14'd1010 : begin out <= 64'b0010101011000010101010001010111000101000110000101010100110100000; end
            14'd1011 : begin out <= 64'b1010011101000010101001010100010000011011010100111010010001000000; end
            14'd1012 : begin out <= 64'b1010010000001010101010100000010100101011101110010010010101111001; end
            14'd1013 : begin out <= 64'b0010011010000110001000100111100010010010110001010010100101011101; end
            14'd1014 : begin out <= 64'b1001111111000111001010011001000110101000000010010010101001110100; end
            14'd1015 : begin out <= 64'b0010011000111011001000000110011010100101110110110010011010000001; end
            14'd1016 : begin out <= 64'b1010100110011011101001010110110010101001011111110010100001110101; end
            14'd1017 : begin out <= 64'b0010000011101111101010011001111110011011010000101010101000101000; end
            14'd1018 : begin out <= 64'b1010101001001100101000000010010110101010000100111010101111100000; end
            14'd1019 : begin out <= 64'b0010100000011101101010111011000100101010110000000010101110111101; end
            14'd1020 : begin out <= 64'b1010101111010100101000101001000100100110101110110010101111000100; end
            14'd1021 : begin out <= 64'b1001100110101101001010110010001000100011001011011010011100011000; end
            14'd1022 : begin out <= 64'b0010100101101101001010110001100110011110110000001010100000101010; end
            14'd1023 : begin out <= 64'b1010000111101000101010000101101000101000111100001010100100110101; end
            14'd1024 : begin out <= 64'b1010101110101001001001111010010110100101011000010010101101010010; end
            14'd1025 : begin out <= 64'b1010000101001111001001100010101010101001100000010010100100101011; end
            14'd1026 : begin out <= 64'b1010110000001110101001001001011100100100111101110010100011011011; end
            14'd1027 : begin out <= 64'b0010011010100010101010100011001000100001011001101001100011000000; end
            14'd1028 : begin out <= 64'b1001111000111110100110101110000010101010101110101010100111001111; end
            14'd1029 : begin out <= 64'b0010010001001010001010000110001010011110000010111010011110000000; end
            14'd1030 : begin out <= 64'b1010000110110000101010010011111000101000111010100001111010011010; end
            14'd1031 : begin out <= 64'b1010100010011011000111100001011010101000111110010010001011010010; end
            14'd1032 : begin out <= 64'b1010000111010010001010000000100000101011010110000010100110100101; end
            14'd1033 : begin out <= 64'b0010101010001100001010101000110010100100010000011001100000001001; end
            14'd1034 : begin out <= 64'b0010100101111011101001111100011010100010110110110010101010000001; end
            14'd1035 : begin out <= 64'b0010010100100000000110011110000010101011100100010010001011001011; end
            14'd1036 : begin out <= 64'b0001000000010010001001011101101100011101000011101001100110011101; end
            14'd1037 : begin out <= 64'b0010001111011000101010101111010010100010011110010010100011010101; end
            14'd1038 : begin out <= 64'b1010101100100100001000100010000110101000101100011010001011100111; end
            14'd1039 : begin out <= 64'b0010010010100100001010111101100110101011101011010001101011001001; end
            14'd1040 : begin out <= 64'b0010010101000010101001011000011110101000001001001010100111101101; end
            14'd1041 : begin out <= 64'b0010010110110110000101000110111100101000111111001010010010010100; end
            14'd1042 : begin out <= 64'b0010000110000010001001000111001000101011010110010010100111110111; end
            14'd1043 : begin out <= 64'b0010100101000001001010001011010000100000010000111010000100110111; end
            14'd1044 : begin out <= 64'b1010100111101100101010110010011000101010110100011001110010100011; end
            14'd1045 : begin out <= 64'b1010101100101111000110100010001010101011111110001010010100000110; end
            14'd1046 : begin out <= 64'b1010101000110011001010111011101100100000101111100010100010011101; end
            14'd1047 : begin out <= 64'b1010101000010100101001000000111100101010000100001010100110101010; end
            14'd1048 : begin out <= 64'b0010001011111101101010011101001010011111110111010010101001110000; end
            14'd1049 : begin out <= 64'b0010100010110101101000000011100010100111110011111001110001001100; end
            14'd1050 : begin out <= 64'b0010100011001100101010101111001010100000010010101010100010000000; end
            14'd1051 : begin out <= 64'b1010010001101001000111000001110010100111110010111010100101011111; end
            14'd1052 : begin out <= 64'b0010101011110010101000001011001000100111000011010010100011100101; end
            14'd1053 : begin out <= 64'b0010100110011000100110111000111110101001001001100010101111101110; end
            14'd1054 : begin out <= 64'b1010011011111011101001111010100100101010110000000010011110000011; end
            14'd1055 : begin out <= 64'b0010011010110110101001011001010000101001010010010010100000111010; end
            14'd1056 : begin out <= 64'b1010001001001000001001101001100100100110101011101010010110100011; end
            14'd1057 : begin out <= 64'b0010101000100100101010100100110010100111010101110010100011010010; end
            14'd1058 : begin out <= 64'b0010101000000110001010100101100110101010111001001010010001110111; end
            14'd1059 : begin out <= 64'b0010100010001111000110001111010110101001011001100010101011010101; end
            14'd1060 : begin out <= 64'b1010100001000100101011000000110000100100111000011010000111111110; end
            14'd1061 : begin out <= 64'b0001000010110001100111001001111000101010011000010001111001110110; end
            14'd1062 : begin out <= 64'b0001100110010001001010001111011010011100000010010010001011001000; end
            14'd1063 : begin out <= 64'b1000111100111001001000000110111000100010110010001010011100110011; end
            14'd1064 : begin out <= 64'b0010100101001011101000001111001110101011101111001010001100000001; end
            14'd1065 : begin out <= 64'b1010101000110001101000110011110100101001100011111001111101010101; end
            14'd1066 : begin out <= 64'b0000010001011101101010110011111010101001010011111010011011111101; end
            14'd1067 : begin out <= 64'b1010100000111000001010100000001000101001100011011001101010011100; end
            14'd1068 : begin out <= 64'b1010100011000010001010000001111010100111101001011010011110001111; end
            14'd1069 : begin out <= 64'b1010101100010011101001001000101100100000000101100010000011110100; end
            14'd1070 : begin out <= 64'b1010100000101011001001111111101010101000011111010001100011001000; end
            14'd1071 : begin out <= 64'b1010101111100011001010101011101010101001000110101010000010011110; end
            14'd1072 : begin out <= 64'b1010101000011011101010101010001010100000111001001010011011110100; end
            14'd1073 : begin out <= 64'b1010100100001111001010111000110100101011111110011010100011101110; end
            14'd1074 : begin out <= 64'b1010010101000110100111100000101110101010100110010010000011110000; end
            14'd1075 : begin out <= 64'b1010100101000000001000001111010100100100010000100010100111111000; end
            14'd1076 : begin out <= 64'b1010101101011111001001001101000100101001010110010010001011000100; end
            14'd1077 : begin out <= 64'b1010100001000011000011110111100110101010100011011010110000001011; end
            14'd1078 : begin out <= 64'b1010100100111111101001101010100010101011101100011010100101011110; end
            14'd1079 : begin out <= 64'b1010001001000000001010101100010010100110000000010010100101101100; end
            14'd1080 : begin out <= 64'b1001101001011100101010010101111110100101001001010010101010000010; end
            14'd1081 : begin out <= 64'b1010001001010001001010110111010110101010110000000010100100100101; end
            14'd1082 : begin out <= 64'b0010100101101000101010010000111100100000011111010010101010110110; end
            14'd1083 : begin out <= 64'b0010011101011010100101101111101110100000000011110010011011101100; end
            14'd1084 : begin out <= 64'b0010101110011010100110100100010110101000001010101001101101011001; end
            14'd1085 : begin out <= 64'b0010101000011111101001011100010110100000000101001010010011010011; end
            14'd1086 : begin out <= 64'b0010011001110010101010000010001100101010111111100010101000001001; end
            14'd1087 : begin out <= 64'b1010011001001010101000111000100010101001000111001010101010001101; end
            14'd1088 : begin out <= 64'b0010101101100011001001111010011110101000111010011010001111110111; end
            14'd1089 : begin out <= 64'b0010011010110000001001100111011110101011110111000010000110000101; end
            14'd1090 : begin out <= 64'b1010011000011111001010100001111010101000001101011010100110111111; end
            14'd1091 : begin out <= 64'b0001001010101111001010001101100010101000110100010010100011001101; end
            14'd1092 : begin out <= 64'b1010100000101001101000100101010110100010100111101001011000111011; end
            14'd1093 : begin out <= 64'b1010100011011001001010110101100010101001000001111010010010111111; end
            14'd1094 : begin out <= 64'b0010101010101010001010010100011110101001110111011010011001100101; end
            14'd1095 : begin out <= 64'b0010101100101101100110010010110100100011100101110010001100111010; end
            14'd1096 : begin out <= 64'b1010101101110001001000010100101110011101000100100010100101001010; end
            14'd1097 : begin out <= 64'b0010010000000010001001010010110000100101101111100001110111000100; end
            14'd1098 : begin out <= 64'b1010101110111011101000110111000100101001000101111010101011110110; end
            14'd1099 : begin out <= 64'b1010000111101110101000101000101000100111111101010010100111001111; end
            14'd1100 : begin out <= 64'b0010100100011010101010011100101110011000001010011010101100100001; end
            14'd1101 : begin out <= 64'b1010101011010010101001101101010100100010101010000010100101010000; end
            14'd1102 : begin out <= 64'b1010001010011000101010010100101010011110111011011010101101011100; end
            14'd1103 : begin out <= 64'b0010100010000101101001011001110100101000100010011010100100011010; end
            14'd1104 : begin out <= 64'b1010100001110000101000010110001010101001001101010010100010011010; end
            14'd1105 : begin out <= 64'b0010101100010111001010011101000100101010011101000001110001001000; end
            14'd1106 : begin out <= 64'b0010100101100000101001001110100100101001100110111010011000110001; end
            14'd1107 : begin out <= 64'b0010100011100000101001000100111010100110100100000010100010110001; end
            14'd1108 : begin out <= 64'b1010001000111011101010001110100000101011110001100010011011110000; end
            14'd1109 : begin out <= 64'b0010100111001010101000000000011010101011010001110010100101000100; end
            14'd1110 : begin out <= 64'b0010100110101001001010100110101110101010011100001010010100111110; end
            14'd1111 : begin out <= 64'b1010010010101010001010010100111010101000000011101010100100110100; end
            14'd1112 : begin out <= 64'b1010011010101011001001011011110110101011111001001010011011111111; end
            14'd1113 : begin out <= 64'b0010011001000011101001010110001110101010001000001010100111111001; end
            14'd1114 : begin out <= 64'b0010100101111110001001100000010010101011111010000010011010011100; end
            14'd1115 : begin out <= 64'b0010011101100011101000000010011100100001000001100010101011111110; end
            14'd1116 : begin out <= 64'b1010000110101011001010010100110000101010000011101010100100011010; end
            14'd1117 : begin out <= 64'b0001100011001100001010110100011010101001010000011010000100100001; end
            14'd1118 : begin out <= 64'b1010100100111011101000000000101010100000110101011010010101000100; end
            14'd1119 : begin out <= 64'b0010000110101101001001011100001110100001111001100010100100011001; end
            14'd1120 : begin out <= 64'b1010100001111010001000001110000100100110110011001010001111001001; end
            14'd1121 : begin out <= 64'b1010101001000000101001110110001110101011011110110010010011100011; end
            14'd1122 : begin out <= 64'b1010100111111101101000000010010110100100000111100001100000011001; end
            14'd1123 : begin out <= 64'b1010011110100101001000010000000110100101111000111010100101110010; end
            14'd1124 : begin out <= 64'b1010000010000100101010011110010010101001010110111010000110100110; end
            14'd1125 : begin out <= 64'b0010101000111011101010001001111010101010100110100010011000111111; end
            14'd1126 : begin out <= 64'b1010101100000011101010000000011100100101001010101010100010101000; end
            14'd1127 : begin out <= 64'b1010011111100100001000110001000110100111101000111010010011111000; end
            14'd1128 : begin out <= 64'b1010100101100100101010010001110110100110110001000010001110101100; end
            14'd1129 : begin out <= 64'b1010010010010100101001001001010100101010001101001010001010110110; end
            14'd1130 : begin out <= 64'b1001100101011001101010101110100010101001100110100010101111011110; end
            14'd1131 : begin out <= 64'b0010100111011001101001100001111100100001101001011010101100101110; end
            14'd1132 : begin out <= 64'b1010001000011010101000000100101100101011111110010010000000000100; end
            14'd1133 : begin out <= 64'b0010100101101100001010011100100100101001011110011010101100011001; end
            14'd1134 : begin out <= 64'b1010101011100100001011000110010010100001000001000010100100001111; end
            14'd1135 : begin out <= 64'b0010010111010110001001111100100110101010000010100010100101001011; end
            14'd1136 : begin out <= 64'b1001110011100100001000001111101010101011010001101010100100011011; end
            14'd1137 : begin out <= 64'b0010101011110110101010110111100010100001100010010010001000101101; end
            14'd1138 : begin out <= 64'b1010100100011101001001101010010000011101101110100010100000100010; end
            14'd1139 : begin out <= 64'b0010100011011011001000110111011010100100010010010010101001111011; end
            14'd1140 : begin out <= 64'b1010101110101111100010101101011010100010110000110010001000011110; end
            14'd1141 : begin out <= 64'b0010101010001011001010010101010110101001111001010010101000100101; end
            14'd1142 : begin out <= 64'b1010101001011101001010101010011010101001000010111010100100000001; end
            14'd1143 : begin out <= 64'b0010100011001100101010000101100100101011010100001010100001011111; end
            14'd1144 : begin out <= 64'b1010100111011110001000001000111010100010011110100010000110011001; end
            14'd1145 : begin out <= 64'b1010011011101011001001100101000010100100011011101010010100011111; end
            14'd1146 : begin out <= 64'b0010101111111001101010110101110010101000010001001010100010110111; end
            14'd1147 : begin out <= 64'b0010101110011110101011000001000110101010111110001010101011000010; end
            14'd1148 : begin out <= 64'b0010100100000011101010011111011010100110100111100001100100000011; end
            14'd1149 : begin out <= 64'b0010101110011111101010100101110100101000100100011010101011101110; end
            14'd1150 : begin out <= 64'b1010100101000000101001011101111000101011100011100010101001101100; end
            14'd1151 : begin out <= 64'b0010101011011010101010011111000100101001010100000010100110001111; end
            14'd1152 : begin out <= 64'b1010100101100111001000010110011010101010001101101010010100010101; end
            14'd1153 : begin out <= 64'b0010100000010011001010000000110010100011100001100010000110001000; end
            14'd1154 : begin out <= 64'b0010011000000110001001111001100010100100110110010010001011111010; end
            14'd1155 : begin out <= 64'b0010001101000110000111101001111010101010011111001010100010101111; end
            14'd1156 : begin out <= 64'b0000001011101111001010110001100000101010100110001010000101011100; end
            14'd1157 : begin out <= 64'b0010101001110111101010010000010100100101100100110010010000011110; end
            14'd1158 : begin out <= 64'b1010011011110000101010001011010100101010000011110010110001000010; end
            14'd1159 : begin out <= 64'b1010010110111101101010010111001010100111010001111010010001001001; end
            14'd1160 : begin out <= 64'b1010101010011011100110101101011100101011010111101010100100101100; end
            14'd1161 : begin out <= 64'b1010011011110010001000110001000000101011010110110010010010000110; end
            14'd1162 : begin out <= 64'b1010101110000101101000001101010100100111100001100010000110010101; end
            14'd1163 : begin out <= 64'b1010101010011110101010000101001100101000101110111010101110101011; end
            14'd1164 : begin out <= 64'b1010101101101001001001101101111110101010010101101010101101011001; end
            14'd1165 : begin out <= 64'b1010100110011000001000110001000000100100011101011010100010101110; end
            14'd1166 : begin out <= 64'b1010011010110011000100100100000000100011011010101010101010000001; end
            14'd1167 : begin out <= 64'b1010100010110001001001110101110000100011011001010001011101010101; end
            14'd1168 : begin out <= 64'b0010100100100000000000110011010000101001110000001010000111101000; end
            14'd1169 : begin out <= 64'b0010101100010010001000001000011110100011010000011010001101011000; end
            14'd1170 : begin out <= 64'b0010100001111010001010100111001110101010000000001010101111111110; end
            14'd1171 : begin out <= 64'b1010100100100001101000100100011100100010111101111010100001101011; end
            14'd1172 : begin out <= 64'b1010100011000001101000001000010010101011100100100001010101010101; end
            14'd1173 : begin out <= 64'b0010011101100110101000001000001110100010101110101010101011100111; end
            14'd1174 : begin out <= 64'b0010101100000001101010111100101010100000001101111010011111111010; end
            14'd1175 : begin out <= 64'b1001111110001101001010000010111110101001110001011001100110111101; end
            14'd1176 : begin out <= 64'b1010100001001010100101010010101000101010011011100010101101100100; end
            14'd1177 : begin out <= 64'b1010010111100010001010100100111100010011010101000010010111100100; end
            14'd1178 : begin out <= 64'b1010010000010010101001110111010000100110000110010010010001000010; end
            14'd1179 : begin out <= 64'b0010100001011111101000101100100010101010000101001010101110100011; end
            14'd1180 : begin out <= 64'b0010101110110100101001001110001000010111000010010010100111101010; end
            14'd1181 : begin out <= 64'b1010001101111000101010100110011100101010110001101010100100100110; end
            14'd1182 : begin out <= 64'b0010001100101011001011000011101010100001111010001010011001010001; end
            14'd1183 : begin out <= 64'b1010001011110001101001011000101110101011110110100001110000001010; end
            14'd1184 : begin out <= 64'b0010011110010101001001000100110110101010111000100010101101001100; end
            14'd1185 : begin out <= 64'b0010101100101011001001010000011100101000010110010010011011010101; end
            14'd1186 : begin out <= 64'b1001111001111101101001001011010000100100110110111010110000001101; end
            14'd1187 : begin out <= 64'b0010101010110101101010101001010010101011101011101010000110010001; end
            14'd1188 : begin out <= 64'b0010000010011010101001000000011000101010001011111010101010111101; end
            14'd1189 : begin out <= 64'b0010100100000110001010100101100010100110011010001010010100011010; end
            14'd1190 : begin out <= 64'b0010000101110001101010010100110100101001001100000010101111010101; end
            14'd1191 : begin out <= 64'b1010001010000000001001000010000100101010000111010010100101110000; end
            14'd1192 : begin out <= 64'b0010101011000001001010101110100010100100011110000010101101000110; end
            14'd1193 : begin out <= 64'b0010101001010100000111111010111000101000100110001010000101001101; end
            14'd1194 : begin out <= 64'b1010100001011111001010001000110010101010000000101010100110110100; end
            14'd1195 : begin out <= 64'b0010011101000110001000101001101110101010100011011010100001101010; end
            14'd1196 : begin out <= 64'b0010010001101000001010100110101100101001011010010010101101101010; end
            14'd1197 : begin out <= 64'b1010010100110011101010011010011100100001110001011010001111000111; end
            14'd1198 : begin out <= 64'b1010011111100000001000101111100110100101111111111010010101010110; end
            14'd1199 : begin out <= 64'b1010101011110111101010010110001010101000000111010001110001110011; end
            14'd1200 : begin out <= 64'b1001111011111001101010101100100010100100100110101010101101010110; end
            14'd1201 : begin out <= 64'b1010101101111101101001101001100000101011101110101010101011001010; end
            14'd1202 : begin out <= 64'b0010100110001101101000111011010000100001010111100010101001101111; end
            14'd1203 : begin out <= 64'b0010101010100000101010100111011000101010001110001010000111100101; end
            14'd1204 : begin out <= 64'b0001110000101110001001010010000000101010101111001010101111111110; end
            14'd1205 : begin out <= 64'b0010100110011000001001100110001110100100011110100001101011000010; end
            14'd1206 : begin out <= 64'b1010100101111110000110101001100000100101011011011010101111001111; end
            14'd1207 : begin out <= 64'b0010101100111000101001001111001100101010111011011010011100101110; end
            14'd1208 : begin out <= 64'b1001110011001001001000110011000100101001101001100010101011010100; end
            14'd1209 : begin out <= 64'b1010000010010011001010110000000110100100101011100010100110110011; end
            14'd1210 : begin out <= 64'b0010100110010101101000010111010110101000011111000010010111011100; end
            14'd1211 : begin out <= 64'b0010100111011111001000101110011010011101000110011010010111101110; end
            14'd1212 : begin out <= 64'b0010101000101101001010001011101000101010111010010010010111101000; end
            14'd1213 : begin out <= 64'b1010100001100111001010010100000110100100001101000010100101111011; end
            14'd1214 : begin out <= 64'b0010011010100010100111010111011010101001000101100010010011001101; end
            14'd1215 : begin out <= 64'b1010001100011100000111101001101100100101000001101010010010110110; end
            14'd1216 : begin out <= 64'b0010010000001000101001110010101100101000000111010010010011001111; end
            14'd1217 : begin out <= 64'b0001110100101100001010001010011110100101001001100010011001001011; end
            14'd1218 : begin out <= 64'b0010101110010101001010110110111010100010000000101010101101001010; end
            14'd1219 : begin out <= 64'b1010001010101100101010100011000110101011100000110010010110011011; end
            14'd1220 : begin out <= 64'b1010011001110001001010000101011000100001001101111010101110001001; end
            14'd1221 : begin out <= 64'b1010100101101001101010110101010100101011010110101010010001010001; end
            14'd1222 : begin out <= 64'b0010101010100000001010001001100110101011110101101010101001010100; end
            14'd1223 : begin out <= 64'b1010101101001011001001101010101100101011100100011010011011100101; end
            14'd1224 : begin out <= 64'b1010100001011110001001000010110100011110110110010010011011011011; end
            14'd1225 : begin out <= 64'b1010010100101111001000001001101110101010010111011010101000111100; end
            14'd1226 : begin out <= 64'b1010100011101001101000001011110110101010111001011010011000010011; end
            14'd1227 : begin out <= 64'b0010010011001011101010100011111100100111110000011010010111001110; end
            14'd1228 : begin out <= 64'b0010011100011000100111111110100110101011111110000001101010100000; end
            14'd1229 : begin out <= 64'b0010010011110000001000001010011010101010001011111010001010111010; end
            14'd1230 : begin out <= 64'b0010100011000010001001111100111110101000010001110010101011110110; end
            14'd1231 : begin out <= 64'b0010011010001000001010110001000110011111111101111010100011101011; end
            14'd1232 : begin out <= 64'b0010101001111001001001000101100010100101100000100010101110001010; end
            14'd1233 : begin out <= 64'b1001110101001010001011000010110000100110010000101010101000101010; end
            14'd1234 : begin out <= 64'b1001111010111100001010101010110000100110100011001010011110001011; end
            14'd1235 : begin out <= 64'b0010011011111000001000110110111100101010011101001010010110000011; end
            14'd1236 : begin out <= 64'b0001110010111000101010001011000000100011000001010010101001011111; end
            14'd1237 : begin out <= 64'b1010101111111100001011000101110010101011100110110010101101000111; end
            14'd1238 : begin out <= 64'b0010100010001001001010111100100000101000101010101010100010011100; end
            14'd1239 : begin out <= 64'b0010010100101110101000111110110100100111100011110001111010010110; end
            14'd1240 : begin out <= 64'b1010100110011010101010100001110000101010101110100010010101001001; end
            14'd1241 : begin out <= 64'b0010100001011001001001000101110110100001011110111010001000001101; end
            14'd1242 : begin out <= 64'b0010101000110101101010111001001110100101000110010010011100010011; end
            14'd1243 : begin out <= 64'b1010100101001011101010110100110000101010111111100010101010000110; end
            14'd1244 : begin out <= 64'b0001111111000100101010101100001010100010011110011010101001001011; end
            14'd1245 : begin out <= 64'b0010011000000101001000010001000110101001110111111001111011100101; end
            14'd1246 : begin out <= 64'b0010101001011000001010000000111000100111001100100010101000001100; end
            14'd1247 : begin out <= 64'b0010110000000100001000010111111010101011101010100010011100101000; end
            14'd1248 : begin out <= 64'b0010011111010110001000000101100100101010101101101001011101001111; end
            14'd1249 : begin out <= 64'b1010001011100000001001101111110100101011010110100010101100101011; end
            14'd1250 : begin out <= 64'b0010101000100111100111100111001000101010000010101010001001100100; end
            14'd1251 : begin out <= 64'b1010101001110011001010101111001000100110110000100001101110011001; end
            14'd1252 : begin out <= 64'b1001001011011001101001100101100000100000111100100010011011000011; end
            14'd1253 : begin out <= 64'b1010100000011101101010100010010010101000110100110010101010101110; end
            14'd1254 : begin out <= 64'b1010100110111001101000000111001000100111010001100010101100110110; end
            14'd1255 : begin out <= 64'b1010001101011011001010111010111110101010111010011010100111000110; end
            14'd1256 : begin out <= 64'b1010101000001001001001000101110000011111011011000010110000000010; end
            14'd1257 : begin out <= 64'b0010101111011101101001010011010110100101111111110010011011101000; end
            14'd1258 : begin out <= 64'b1010100010111110001010100100101110011100101011101010101010001010; end
            14'd1259 : begin out <= 64'b1010100100010011001010100101001010011101101110000010100100010011; end
            14'd1260 : begin out <= 64'b1010101001011010101000000011010110101001110000010010000101000111; end
            14'd1261 : begin out <= 64'b1010100100010010101001100010010010101011110100110010101000001000; end
            14'd1262 : begin out <= 64'b0010011100000101101010000001100010101000100100100010101001011110; end
            14'd1263 : begin out <= 64'b0010001010010110101010001010001110100101100011001010100100101100; end
            14'd1264 : begin out <= 64'b1010010000110110101010111010011100101000000000101010101101011110; end
            14'd1265 : begin out <= 64'b1010000000111001101010001101000100101001111011001010000110101100; end
            14'd1266 : begin out <= 64'b1010110000011001101001100101010110101011011100001010010001111101; end
            14'd1267 : begin out <= 64'b0010011011111011001001100111110110101010001001101010001110100110; end
            14'd1268 : begin out <= 64'b1010100011000011101010011101001010101010100111101010100101100000; end
            14'd1269 : begin out <= 64'b1010011110101010101010010010001100011001110001100010000100011000; end
            14'd1270 : begin out <= 64'b0010011110000001101010010111010010100111001001110010011111100110; end
            14'd1271 : begin out <= 64'b1010101010101000101001100100000110101000000111100010010110000100; end
            14'd1272 : begin out <= 64'b0000000110011000000111101001111010011001010100111010010101010100; end
            14'd1273 : begin out <= 64'b1010101100001110101010011100001100100100110010110001100101010011; end
            14'd1274 : begin out <= 64'b0010000010101101101010011011100100101000001110010010101101101001; end
            14'd1275 : begin out <= 64'b0010010111110010101010110001111010010111111111000010000110101100; end
            14'd1276 : begin out <= 64'b1010100000111100101010100011011100100011001010001010010110011100; end
            14'd1277 : begin out <= 64'b0001100010111010001010110000011100101011001110111010100010110000; end
            14'd1278 : begin out <= 64'b1010010000111000101010011010110100011100101010100010100010110110; end
            14'd1279 : begin out <= 64'b0010101100100111101010010111101000101010011010100010100011001101; end
            14'd1280 : begin out <= 64'b0010100010101100101010110000001010100101101110100010000111111001; end
            14'd1281 : begin out <= 64'b0010000111110000101010100010110100100111100011100010010100001001; end
            14'd1282 : begin out <= 64'b0010010100010111101010111110110010101001110011011010001100011000; end
            14'd1283 : begin out <= 64'b1001110111011100101001110100101110101000011111111010100111001000; end
            14'd1284 : begin out <= 64'b0010101110011010101001000001101110101000011010011010101100011001; end
            14'd1285 : begin out <= 64'b1010100111011101001000100010110000100100111111111010100101111011; end
            14'd1286 : begin out <= 64'b1010100111001101101010000001001010100111010100011010101100001001; end
            14'd1287 : begin out <= 64'b1010000111001100001010100100101100100010000101111010100100000011; end
            14'd1288 : begin out <= 64'b1010000010101010001010010100101000100101000001100010011010000010; end
            14'd1289 : begin out <= 64'b0010101100001011101010001101110110100100010011000010100111001101; end
            14'd1290 : begin out <= 64'b1010110000001101001010110010111100011010001101011010101000111100; end
            14'd1291 : begin out <= 64'b0010100010100011101010010100001100101001000110111010001000001000; end
            14'd1292 : begin out <= 64'b0010010101001000001000111101001100101010011000000010000011010100; end
            14'd1293 : begin out <= 64'b1010100001111001001000011001110000101000011001111010010101000110; end
            14'd1294 : begin out <= 64'b0010100100010111101001011100010000101010100011101010010101011110; end
            14'd1295 : begin out <= 64'b1010011100011010101000000101001100101010000010100010010011110110; end
            14'd1296 : begin out <= 64'b1010101101000000001010001010111010100101110000110010100000000111; end
            14'd1297 : begin out <= 64'b1001111000001011101000110000010100100101010101101010001011110111; end
            14'd1298 : begin out <= 64'b1010010110001010101010011110011010101011101011110010101111000111; end
            14'd1299 : begin out <= 64'b1010011000110000001010000001000110101001100100001010011100110000; end
            14'd1300 : begin out <= 64'b1010011110111100001010000001111110100110010011110010101111111010; end
            14'd1301 : begin out <= 64'b1010001111000000001010101110011000101001010001100010100001111010; end
            14'd1302 : begin out <= 64'b0010101011111000001010010011000000100111110001001010101010100100; end
            14'd1303 : begin out <= 64'b1010101111011111001001011010011110101001101110000010100010001110; end
            14'd1304 : begin out <= 64'b1010100110011100100111010100011010100110001011100010010110001101; end
            14'd1305 : begin out <= 64'b1010100110100001001010101010001000101000100101000001111101111101; end
            14'd1306 : begin out <= 64'b0010100111010111000111011101011110011101101101001010101101100010; end
            14'd1307 : begin out <= 64'b0010000110100111100101000011111110010111111010011010101010110101; end
            14'd1308 : begin out <= 64'b1010100000110010001010111111011100101000010110100010010100011011; end
            14'd1309 : begin out <= 64'b1010101011101001101010111110110000101001010110011010011110111001; end
            14'd1310 : begin out <= 64'b1010001011101001001001001100010100101000001100111010011101011010; end
            14'd1311 : begin out <= 64'b0010010010111010101010111010110100100110100101101010001100001011; end
            14'd1312 : begin out <= 64'b1010101111001100001001111000110110100111011110000010101000000101; end
            14'd1313 : begin out <= 64'b0010010111010000101010001000001110100010111000110000110011100100; end
            14'd1314 : begin out <= 64'b0010101110111101101010111100111010101000101100100010011001010111; end
            14'd1315 : begin out <= 64'b1010101010110001101010011100110110101000100111000010101101001011; end
            14'd1316 : begin out <= 64'b1010100010111010001010100111001100101011101110001010101111111000; end
            14'd1317 : begin out <= 64'b1010010001000010101010101110000100100111110010110010100110100000; end
            14'd1318 : begin out <= 64'b0010011010101001101001101111000110100110011111100010100101010010; end
            14'd1319 : begin out <= 64'b0010100100000110001010011110001100011111001000011001111010100111; end
            14'd1320 : begin out <= 64'b1010101100000010001010010110010100101011010100000010101011110001; end
            14'd1321 : begin out <= 64'b0010000100001110001010101011000110101001111100110010101110011001; end
            14'd1322 : begin out <= 64'b0010100010001100101010011110111100100110001001111010101000011111; end
            14'd1323 : begin out <= 64'b1010101111010101101010110000101000100000010111110001101101100101; end
            14'd1324 : begin out <= 64'b1010101100101010001001010000000000101011111101011010100111001100; end
            14'd1325 : begin out <= 64'b1010101111010101001010001100001100100100011001001010101101010100; end
            14'd1326 : begin out <= 64'b1001101000100011100110010100111010100101000010110010011111001100; end
            14'd1327 : begin out <= 64'b1010000001110101101010101001111000011001110111111010010001011100; end
            14'd1328 : begin out <= 64'b0001110100010000001001110010101010101000101110111010101110100100; end
            14'd1329 : begin out <= 64'b0010001110100011001010110001111100100100101001110010101010011011; end
            14'd1330 : begin out <= 64'b0010001101101011001010100010011110100011110010001010101000011110; end
            14'd1331 : begin out <= 64'b0010011100010101001000110101110110101010110000101010000101010101; end
            14'd1332 : begin out <= 64'b0010101010111101001010110010010100100001111100100010100011010100; end
            14'd1333 : begin out <= 64'b0010100000111000101001011110100010100000011100000001011011101010; end
            14'd1334 : begin out <= 64'b1010101001011011101001010000101100101011001111101010100000111101; end
            14'd1335 : begin out <= 64'b1010100000011011001010100001010000101000000010011010001111100010; end
            14'd1336 : begin out <= 64'b1001110110110110101010011110000100101011101110011010101011101110; end
            14'd1337 : begin out <= 64'b1001100100101101101001111000010010100111000011100010011100000101; end
            14'd1338 : begin out <= 64'b0010101011110000101001000010110010101001111100001010101001111111; end
            14'd1339 : begin out <= 64'b1000101100010111001001111111011100011010110110000010010001100100; end
            14'd1340 : begin out <= 64'b0010001010000111001010010111100100011011101111000010010111100000; end
            14'd1341 : begin out <= 64'b0010010010100110001001011011101100101000110001111010100001010111; end
            14'd1342 : begin out <= 64'b1010011010010100101001010101101110101011101100100010011111010111; end
            14'd1343 : begin out <= 64'b0010100101010111101010110011110100101001111100100001110110101110; end
            14'd1344 : begin out <= 64'b1010101101101001001000011001010010101010101001101010011000100100; end
            14'd1345 : begin out <= 64'b1010010011001001001010101010011010101000100000100010101010111001; end
            14'd1346 : begin out <= 64'b1010101001000011101010100000000000100110101000110010001000110000; end
            14'd1347 : begin out <= 64'b0010100000000011001001110000101000101001000111111001101110100010; end
            14'd1348 : begin out <= 64'b1010000010001101101010010010101010100011010111000010001110100001; end
            14'd1349 : begin out <= 64'b1010101011010110101001111010110010101000111001011010101101110110; end
            14'd1350 : begin out <= 64'b1010011010011111001010110011000010100101000111010010010110000010; end
            14'd1351 : begin out <= 64'b0001010100100100100110100000111010101011101110010010000010001010; end
            14'd1352 : begin out <= 64'b0001000101110100101010111011000110101001101001110010011101010011; end
            14'd1353 : begin out <= 64'b0010000100100010101001011011111010011101001010110010101000001010; end
            14'd1354 : begin out <= 64'b0010000101101110101001011101111010100110100100001010101110100001; end
            14'd1355 : begin out <= 64'b1010100001001010101010100010010100101011001110010010101000110001; end
            14'd1356 : begin out <= 64'b0010101000110000101010000001111000101011111110001010010111110000; end
            14'd1357 : begin out <= 64'b1010011100111101101000110100000110101000101111010010011000101010; end
            14'd1358 : begin out <= 64'b1010101000010001101000110100110110101010010111100010000001000001; end
            14'd1359 : begin out <= 64'b0010101111111000101010000110111110100100010101010010000111110101; end
            14'd1360 : begin out <= 64'b0010100011101000001001111111100010101011001000111010001001110100; end
            14'd1361 : begin out <= 64'b1010011111001101001010100100010010101000001010101001101010111011; end
            14'd1362 : begin out <= 64'b0010101011000000000110101011111000101001010100010010001000110101; end
            14'd1363 : begin out <= 64'b1010100101000111001010000010011010100110010100010010001010001100; end
            14'd1364 : begin out <= 64'b0010001000010110001010110011011110101001101101000010101110101000; end
            14'd1365 : begin out <= 64'b0010100011000011001001011011000110011110100110100010010100000110; end
            14'd1366 : begin out <= 64'b0010010010001111001001110010110100100000000000000010010000100110; end
            14'd1367 : begin out <= 64'b1010100001111000101001010111010110101011000100100010101111000001; end
            14'd1368 : begin out <= 64'b1010001111000010000110101110000010101011101100110001001101111111; end
            14'd1369 : begin out <= 64'b1010101011001111001010111101001100011111010001110010010011110010; end
            14'd1370 : begin out <= 64'b1001111001111100001001111011110110100000010111001010000100111001; end
            14'd1371 : begin out <= 64'b1010101011011000101010100000011110100000010010111010100001100100; end
            14'd1372 : begin out <= 64'b1010101001111000001010110111111100001100110110011010010111110000; end
            14'd1373 : begin out <= 64'b1010100110110111001010100010010110100100111100001010101011110011; end
            14'd1374 : begin out <= 64'b0010101010101110101000010011110010101010011110000010010010101001; end
            14'd1375 : begin out <= 64'b1010011000100110101000111001010110101100010110000010100010000111; end
            14'd1376 : begin out <= 64'b0010001000110100001001010011010000100000011001100010001101000010; end
            14'd1377 : begin out <= 64'b0010100111000011001010100001110110100100100011111010100011000011; end
            14'd1378 : begin out <= 64'b1010100000111101001010010011100000101011101101101010000111100011; end
            14'd1379 : begin out <= 64'b1010010111101101101000111000001000100100101101011001110110000111; end
            14'd1380 : begin out <= 64'b1010011001000101100101001101001110010011110011111010101100000011; end
            14'd1381 : begin out <= 64'b0010011010110101100111001000100010100111110111011010100000001110; end
            14'd1382 : begin out <= 64'b1010011001010111001000100100000000101001110110101010011100000001; end
            14'd1383 : begin out <= 64'b0010100100000011001000010000110110101010010001111010101101110111; end
            14'd1384 : begin out <= 64'b0010101010110110101001111100111000100001011001100010011101110011; end
            14'd1385 : begin out <= 64'b0010100001001100101010011011100010100111110000110010011100100000; end
            14'd1386 : begin out <= 64'b1010101110001101101001110001110110101010110011101010011001010110; end
            14'd1387 : begin out <= 64'b1001010011111110001001011110001110101010001101110010101110110000; end
            14'd1388 : begin out <= 64'b1010101010100001100110100001110000100100000010101010010001100111; end
            14'd1389 : begin out <= 64'b0010011011001011001010110010000010100101011110110010011110101110; end
            14'd1390 : begin out <= 64'b1010000101100100001010001100101000100110010111110010100000001000; end
            14'd1391 : begin out <= 64'b0010101001000111001001111101010000100111111100110010011011000110; end
            14'd1392 : begin out <= 64'b1010101110011001001010011100011000101001101010111010010100001101; end
            14'd1393 : begin out <= 64'b1010010000011001101001010010000010100001001110010010100111100000; end
            14'd1394 : begin out <= 64'b0001111101010001001010110100000100100101100110100010101110111000; end
            14'd1395 : begin out <= 64'b1010011001011001001010110001110010101010010000101010011111011111; end
            14'd1396 : begin out <= 64'b0010100101000101001010010011001000011011001101100010001100110011; end
            14'd1397 : begin out <= 64'b1010100011001110101010000100011010100111011101110010100111001110; end
            14'd1398 : begin out <= 64'b1010100000111011101001010101001000100101011000001010101110011100; end
            14'd1399 : begin out <= 64'b0010100111000001001010011000000000101100001110100010100010101100; end
            14'd1400 : begin out <= 64'b0010101101110001101010101010110100101000011011100010000100100001; end
            14'd1401 : begin out <= 64'b1010101000100100001010100110011010101001111100101001110010010101; end
            14'd1402 : begin out <= 64'b1001011101111000101010110001110000100101011101111010010101111011; end
            14'd1403 : begin out <= 64'b1010100101100110101010110000000000101011011100000010100000010001; end
            14'd1404 : begin out <= 64'b1001010001010111101010100000001010100101000010111010101011110100; end
            14'd1405 : begin out <= 64'b1010101001000001001001001110010100011110001100001010101101111010; end
            14'd1406 : begin out <= 64'b1010010001111001101010101101011100101001000100011010101111110000; end
            14'd1407 : begin out <= 64'b0010100111010001000111111111000100101001111000100010011100100100; end
            14'd1408 : begin out <= 64'b0010101110000001101010000111000000011110000010101010100001100110; end
            14'd1409 : begin out <= 64'b0010011100100111001000011100100000100001011100110010010110011011; end
            14'd1410 : begin out <= 64'b0010101001000111001001101011111110101000011001010010101001000100; end
            14'd1411 : begin out <= 64'b0010010100001001001010000000100100101011111100101010010111011011; end
            14'd1412 : begin out <= 64'b1010100100110111101010111101011110101100000001011010101010110101; end
            14'd1413 : begin out <= 64'b1001100111000010101010111110110100101001110100010010100000000110; end
            14'd1414 : begin out <= 64'b1001110101011001001010011001111100101010011111111001110101100010; end
            14'd1415 : begin out <= 64'b1001110000001101101001000111100010100101011011011010010100111110; end
            14'd1416 : begin out <= 64'b0001100110010111101001111101110110010110110111100001101010101000; end
            14'd1417 : begin out <= 64'b1010101100001000101010110100010100100101000010100010101011010101; end
            14'd1418 : begin out <= 64'b0010001100010001001010110001111110100001101110111010100000101101; end
            14'd1419 : begin out <= 64'b1010101111001111000111110100110010100111001011101010101010011111; end
            14'd1420 : begin out <= 64'b0010101001100001101001111010111110100101001101111010100011001010; end
            14'd1421 : begin out <= 64'b0010101110110100100111001101111100100011011001011010000011010010; end
            14'd1422 : begin out <= 64'b1010001011100100001010101000101000100000101010001010011100101100; end
            14'd1423 : begin out <= 64'b1010101101011010001001101001100000100100011101010010100110101110; end
            14'd1424 : begin out <= 64'b0010000111001101101001111010001110101010110100101010010010101101; end
            14'd1425 : begin out <= 64'b0001101010011100101001110111100000011111100011001010101010010001; end
            14'd1426 : begin out <= 64'b1010000001011111101010001111000110101010101101010010001101100010; end
            14'd1427 : begin out <= 64'b0010101001001101001010100011011110100110110100101010100000010100; end
            14'd1428 : begin out <= 64'b0010011000101110101010101110001100101000011110111001110100110011; end
            14'd1429 : begin out <= 64'b0010010010000001001001110000100100011011001111100010101001101010; end
            14'd1430 : begin out <= 64'b0010100101100000101010101010010010100100000000101010010110100010; end
            14'd1431 : begin out <= 64'b1010100011101100101001101000001110100011011000000010011110111100; end
            14'd1432 : begin out <= 64'b1010100000000011101000111001111010101000100101111010001000001100; end
            14'd1433 : begin out <= 64'b1001111001001010001010011011001100101001000011101010100001111111; end
            14'd1434 : begin out <= 64'b1010011100111011001010100000001000100101011010110010010000111010; end
            14'd1435 : begin out <= 64'b0001111011010000100111000101100110101001001010111010011111100000; end
            14'd1436 : begin out <= 64'b0010101100111110001010000111101000100000000110001010100000001101; end
            14'd1437 : begin out <= 64'b1010101001000011001010001011011100101011110110011010100011000010; end
            14'd1438 : begin out <= 64'b1010010101010010001010101010110000101010111010110010010110001110; end
            14'd1439 : begin out <= 64'b1010100000110001001010010100011100011010101111010001000110001111; end
            14'd1440 : begin out <= 64'b0010000111110100001000101101111000101001011000100010000000100001; end
            14'd1441 : begin out <= 64'b1010000001100111001010001010110000101011111100000010010100111010; end
            14'd1442 : begin out <= 64'b1010100001000010001010010000000100101000100000111001111110010110; end
            14'd1443 : begin out <= 64'b0010100000110100101010110010001100101001010011111001111101111001; end
            14'd1444 : begin out <= 64'b1010101011110100101010111011101100011110010111010001110111001100; end
            14'd1445 : begin out <= 64'b0010000101101110001000000010100000101000000001011010101010100101; end
            14'd1446 : begin out <= 64'b0010010110110000101001111100011010100110101111001010011011000011; end
            14'd1447 : begin out <= 64'b0010100100111010101010001110000010101001010001011010100010110100; end
            14'd1448 : begin out <= 64'b1010001111111000001010001101101100101000101111011010101110100000; end
            14'd1449 : begin out <= 64'b0010010000000011001001001100100010100101011011010010101010101010; end
            14'd1450 : begin out <= 64'b0010101001010101001010001101010000101000110000101010101111111000; end
            14'd1451 : begin out <= 64'b0010011000010011101010010011010100101011011000101010010111011100; end
            14'd1452 : begin out <= 64'b0010100001100101001001001111001110100010110110111010101110110011; end
            14'd1453 : begin out <= 64'b1010010000101011101010110111110100011000101111111010010111011010; end
            14'd1454 : begin out <= 64'b1010011001000010001001010100010100011100110110001010101001001110; end
            14'd1455 : begin out <= 64'b0010011110001101101010000001110100100111001111000010100111101110; end
            14'd1456 : begin out <= 64'b0010000111010101101001011110001100101011011111111010100001010010; end
            14'd1457 : begin out <= 64'b1010010010011000000111011110111110101001000011000010101100100110; end
            14'd1458 : begin out <= 64'b0010100011001010001010111100100110100111000110001001101111101010; end
            14'd1459 : begin out <= 64'b0010100101110110001000100011110010101100000000100000101011101001; end
            14'd1460 : begin out <= 64'b1010100000101010001010100110110010100000111110100010100100110110; end
            14'd1461 : begin out <= 64'b0010101001111011101000001010110000100100101001101010011000010110; end
            14'd1462 : begin out <= 64'b1010101111101101101010100111100010100011111100110010011001000011; end
            14'd1463 : begin out <= 64'b0010101110010001101010111000001110100100100011000010100110000011; end
            14'd1464 : begin out <= 64'b0010011100100111001000010111010000011100000101101010100000101010; end
            14'd1465 : begin out <= 64'b0010101001001101001001000000111110101001001111110010001110000001; end
            14'd1466 : begin out <= 64'b0010101100011011101001001110111000100011101111111001101101000101; end
            14'd1467 : begin out <= 64'b1010010110101010001001011110100110101000000001011010011011011101; end
            14'd1468 : begin out <= 64'b0010101100010101001001011000100000101001111010000010100001100010; end
            14'd1469 : begin out <= 64'b1010101101011111101001011011001010101010010011010010001101010110; end
            14'd1470 : begin out <= 64'b1001110011100101101010110101011100101010110111010010010011111001; end
            14'd1471 : begin out <= 64'b1001111001010111101010011101110100100101011100011010010010011010; end
            14'd1472 : begin out <= 64'b1001101110000001001001110100101010100100100011100010001101111011; end
            14'd1473 : begin out <= 64'b1010100000010011101000010100000100100000011001101010000010100001; end
            14'd1474 : begin out <= 64'b0010010000001001101001111110001100100111011011100010100001000001; end
            14'd1475 : begin out <= 64'b0010101110101010001001100110001000101001110110101010101011111101; end
            14'd1476 : begin out <= 64'b0010010010000010101010000110011000101011000110110010001011111110; end
            14'd1477 : begin out <= 64'b1010101101101111001001001000110100101000110110100001110111110011; end
            14'd1478 : begin out <= 64'b0010100010001101001000000110001000100110111000111001110001101000; end
            14'd1479 : begin out <= 64'b0010101001010001101001010101110000100010110100101010101111010011; end
            14'd1480 : begin out <= 64'b1010100100011111101010100110111110101010111001110010101001110111; end
            14'd1481 : begin out <= 64'b0010100101110101001010000100011100100010111000011010011001010101; end
            14'd1482 : begin out <= 64'b0010100111000100001010011001101000100101110011011010100001010111; end
            14'd1483 : begin out <= 64'b0010010011001011001010011100101000101000110000110010101110010111; end
            14'd1484 : begin out <= 64'b0010001110010010101001000001110100100111111110000010000111010010; end
            14'd1485 : begin out <= 64'b1010010011110000101010011100011100100110011100110010011110100100; end
            14'd1486 : begin out <= 64'b0010011000010101101010111111001010101001111010001010101001101010; end
            14'd1487 : begin out <= 64'b1010101100000111001001111000000100100001010001110001110100010010; end
            14'd1488 : begin out <= 64'b0010000011001000101001001011010010100011111010010001011110111111; end
            14'd1489 : begin out <= 64'b0010101010010100101000101101001010100110100100011010101111010000; end
            14'd1490 : begin out <= 64'b0010100000111010001010111011001000100011001001111010011111100010; end
            14'd1491 : begin out <= 64'b1010100111010111001010001101010100100001000110000000100011010011; end
            14'd1492 : begin out <= 64'b0010010110010011101001011001101100101011110011011010101110101010; end
            14'd1493 : begin out <= 64'b0010101011110110101010001110100010101010100010000001010000010010; end
            14'd1494 : begin out <= 64'b0010100001111011001001111011111110101000000100110010011101001010; end
            14'd1495 : begin out <= 64'b0010101010010110001000101101010110101001011100111010011001000001; end
            14'd1496 : begin out <= 64'b1010101111000011101010011111001100100000001010011010100111100000; end
            14'd1497 : begin out <= 64'b1010001100011011000101100101111010100111010111100010101101100001; end
            14'd1498 : begin out <= 64'b1010100111000000001010100010100100011100111010100010100110100010; end
            14'd1499 : begin out <= 64'b1010011101101011001001100010011110100101101110001010101010011110; end
            14'd1500 : begin out <= 64'b1010101111101001001010111101001110100110010110001010010010110110; end
            14'd1501 : begin out <= 64'b1010101111000101001010000111101010101000101110010010011110010001; end
            14'd1502 : begin out <= 64'b1010010010100111001010101011111010001010111001010010101001101101; end
            14'd1503 : begin out <= 64'b0001111010011011001001100101100000100001100100010010100101010111; end
            14'd1504 : begin out <= 64'b0010010000111111101010000101100000101010101001011010100011111000; end
            14'd1505 : begin out <= 64'b1010100100000010001010110110001110011100000010111010001001001111; end
            14'd1506 : begin out <= 64'b0001111101001000000100001010110110101010100111101010100111001111; end
            14'd1507 : begin out <= 64'b0001111100001001001001100001100110101010001001000010100000101101; end
            14'd1508 : begin out <= 64'b0010100111110110101010111011110010101000100010000010100000111101; end
            14'd1509 : begin out <= 64'b0001100001111110101001110100001000100100001011101001101101111100; end
            14'd1510 : begin out <= 64'b0010100101010010101000000001100000101001001101101010101101100011; end
            14'd1511 : begin out <= 64'b1010100010111001101000100111110000101001011001100010001010011101; end
            14'd1512 : begin out <= 64'b1010100000001110000000101100011110100110110100010001010010111110; end
            14'd1513 : begin out <= 64'b1010101001001010101001010001001100100000101111000010011101110101; end
            14'd1514 : begin out <= 64'b1010100111110011001001011100101000100000101100111001011111010100; end
            14'd1515 : begin out <= 64'b1010010000101010001010011111001100101010110010111010100111001011; end
            14'd1516 : begin out <= 64'b0010010001011000100101011100010010101001011100110010100100011000; end
            14'd1517 : begin out <= 64'b0010100001000111001010100010000010101011110001111010010101111001; end
            14'd1518 : begin out <= 64'b1010010010000100101010101010011110100011110110110010011111001100; end
            14'd1519 : begin out <= 64'b1010100000101111001010010001101010101000011011000001110010000000; end
            14'd1520 : begin out <= 64'b1010101101110101001010110010111110101010010011101010100011111001; end
            14'd1521 : begin out <= 64'b1010100101001100001010101001111010100000100001101010011000100110; end
            14'd1522 : begin out <= 64'b1010101010010110101000111001011000100100011011001010011010100111; end
            14'd1523 : begin out <= 64'b1010101010010001101001111110110100100100011110111010000000010100; end
            14'd1524 : begin out <= 64'b1010100101001111101010110101010000011100000100011010101100010010; end
            14'd1525 : begin out <= 64'b1010101111011000000110101111010100100100111001001001110110110100; end
            14'd1526 : begin out <= 64'b1010100111100101001010000100001110101010101111001010011111110111; end
            14'd1527 : begin out <= 64'b1010101010000110001010010001010010101000001001110010010100100100; end
            14'd1528 : begin out <= 64'b1010100101001100001001010000111100100001011000111001010011101010; end
            14'd1529 : begin out <= 64'b1010101000110000101001100111110000101010000001101010010001110110; end
            14'd1530 : begin out <= 64'b0010101000101111101001001000011100100100111011101010001111110001; end
            14'd1531 : begin out <= 64'b1001111110100000001010110001010010101001001110010001110100000111; end
            14'd1532 : begin out <= 64'b1010101101100100101010111111101100100101001010101010100101111111; end
            14'd1533 : begin out <= 64'b0010011101011111001010010011010110100111110000111010011001110011; end
            14'd1534 : begin out <= 64'b0010100001000011101010110000111000100111000000000010101110100101; end
            14'd1535 : begin out <= 64'b1010101110101110101010001101000010101010010110001010001100000101; end
            14'd1536 : begin out <= 64'b0010010011011110101010011011101100101010110111110010100011010100; end
            14'd1537 : begin out <= 64'b0010100110110001101010111110000110100010001010110010011100011010; end
            14'd1538 : begin out <= 64'b1001110000101001101010010000111010101000001010101010101100110011; end
            14'd1539 : begin out <= 64'b1001110001110000101001010011110000100111000001100010110001100010; end
            14'd1540 : begin out <= 64'b0010101100000010001010011000110100100101011001101010100101101100; end
            14'd1541 : begin out <= 64'b1010101010010110001001101000110010100011001111110010101000001101; end
            14'd1542 : begin out <= 64'b0010101000011100101010011101000000100101101011011010000001110010; end
            14'd1543 : begin out <= 64'b0010011000101001101010100101111000101011011000000010101001100110; end
            14'd1544 : begin out <= 64'b1010100001010011101010101010010000011110100100100010100010000000; end
            14'd1545 : begin out <= 64'b1010101111110010001001111101011000101000101101111010100100110011; end
            14'd1546 : begin out <= 64'b0001110101000010001001110011001100101010110100011010001000010110; end
            14'd1547 : begin out <= 64'b0010100011110111101010111101000100101011010001101010101010011100; end
            14'd1548 : begin out <= 64'b1010001111010100001010000001000100101000011101110001101000100010; end
            14'd1549 : begin out <= 64'b0010010000011110101010100101101110011110101010110010011011110011; end
            14'd1550 : begin out <= 64'b0010101001101011101000000100010110011001110001100010101011011111; end
            14'd1551 : begin out <= 64'b1010101100100101101001101101111000101010100100101010100100100110; end
            14'd1552 : begin out <= 64'b0001110001110100001010010000000100011100100100100010001100111111; end
            14'd1553 : begin out <= 64'b1001011110011100101001111011001010100001111010011010011010001000; end
            14'd1554 : begin out <= 64'b1010100001111001101010000111100110101010100011101010001100100100; end
            14'd1555 : begin out <= 64'b1001111110000010101001011000111100100100011110001010100011100110; end
            14'd1556 : begin out <= 64'b0010100011011011100101110011111110101000001101001010010000100000; end
            14'd1557 : begin out <= 64'b1010101010110000101001101101110000001110011010000010100111110011; end
            14'd1558 : begin out <= 64'b0010100000110000001001110011010010101000011000011010100011101111; end
            14'd1559 : begin out <= 64'b1010101001111000001001100110011010100100011100100010101100110000; end
            14'd1560 : begin out <= 64'b1010101101001000001001101101101110101001101010010010100101001100; end
            14'd1561 : begin out <= 64'b1010011000001001001001011000101110100110111110100010011111010011; end
            14'd1562 : begin out <= 64'b0010100010011101001010000110011000100100011000010010100101111011; end
            14'd1563 : begin out <= 64'b0010101110111100101001100000011100101010100001010010101100000100; end
            14'd1564 : begin out <= 64'b0010011010110001000110111010110010101001101011011010010100010001; end
            14'd1565 : begin out <= 64'b1010101100110011001010010000100010100111010101110010000100001110; end
            14'd1566 : begin out <= 64'b0010101000110101001010010111110000100000110010100010010111101011; end
            14'd1567 : begin out <= 64'b1010100100111111101000100010011010101010000011001010101110000101; end
            14'd1568 : begin out <= 64'b0010000000000010000110111000000110101000110100000010010100101001; end
            14'd1569 : begin out <= 64'b1010011011100010001000100101100100101011011111100010001000010001; end
            14'd1570 : begin out <= 64'b1010100100101111001000110000110110101011000100001001111111100110; end
            14'd1571 : begin out <= 64'b0001100001111100000110000110010100101010111110001010100001110010; end
            14'd1572 : begin out <= 64'b0010000011100010101000011010011100011110000100010010011000111011; end
            14'd1573 : begin out <= 64'b1010011100110101101010001010001000100110001000111010100001100111; end
            14'd1574 : begin out <= 64'b0010000111001000001001101001001000100010000010100010011000001101; end
            14'd1575 : begin out <= 64'b1010011101110100000110101000001110101010000001100010100010001111; end
            14'd1576 : begin out <= 64'b1010101001000100000111111011111010101010111110111001100100001011; end
            14'd1577 : begin out <= 64'b1010101010000011101010011011011000100111001011100010101000000100; end
            14'd1578 : begin out <= 64'b0010100110100001001000000001111100100111011101000010011010000101; end
            14'd1579 : begin out <= 64'b1010101101011000001001101000001000101011000010011010100010100001; end
            14'd1580 : begin out <= 64'b1010100011111011001001000101010010100000101100110010010110001000; end
            14'd1581 : begin out <= 64'b1010010100000010001001110111100110011111111011110010100100101100; end
            14'd1582 : begin out <= 64'b1010101110011000001011000001110110101011001100101010100001000000; end
            14'd1583 : begin out <= 64'b0010101010000000101010001100011110101010011001011010001100000000; end
            14'd1584 : begin out <= 64'b0010100000011111001000000001110000101001000110101010101000010111; end
            14'd1585 : begin out <= 64'b0010100111010101001000010010001100100101000011101010010001011100; end
            14'd1586 : begin out <= 64'b1010010110001101101010101010001110100011001100101010101010000110; end
            14'd1587 : begin out <= 64'b1010010101011010001010010010011000101001000100001010100111010000; end
            14'd1588 : begin out <= 64'b1010011011111111101010001100010110100101111000111010000010111000; end
            14'd1589 : begin out <= 64'b0010011010010100101010001010111100100101101000010001111001000001; end
            14'd1590 : begin out <= 64'b1010011010110110001000110010001010101000100100010010100100101001; end
            14'd1591 : begin out <= 64'b0010100010011110001010100000111110100000000011011010000000110101; end
            14'd1592 : begin out <= 64'b0010011000110101001010011111101100100111110000001010100010000111; end
            14'd1593 : begin out <= 64'b1010100001010010000111000011000010101000101011111010001111101100; end
            14'd1594 : begin out <= 64'b0010101110010011101010110101111010100101000010101010011010001101; end
            14'd1595 : begin out <= 64'b0010101101101011101010100110100110100110001001111010010110011101; end
            14'd1596 : begin out <= 64'b0010011110111000101010001010111110101000010000000010101000001100; end
            14'd1597 : begin out <= 64'b0010000100111001101010011101101110101011101011100010000001101010; end
            14'd1598 : begin out <= 64'b1010100011000110101000010101000110100111001011100010100011010010; end
            14'd1599 : begin out <= 64'b1000111101101100001010101101111010100101001011101010100001101010; end
            14'd1600 : begin out <= 64'b0010101101110010101000110011110100100100010010101010101010010100; end
            14'd1601 : begin out <= 64'b0010011100100000001011000100110110100110101100111001110111011001; end
            14'd1602 : begin out <= 64'b0010101000111111000110100000111000100100111101001010101010001111; end
            14'd1603 : begin out <= 64'b0010100000001000101010110001000000100001000111110010100100111100; end
            14'd1604 : begin out <= 64'b0001100111100101100110011110001100101001110111111010010010000000; end
            14'd1605 : begin out <= 64'b1010001111111101000111010100100110100111101011000010010011011010; end
            14'd1606 : begin out <= 64'b1010011110011100101000110000110010101010111000110001111001001101; end
            14'd1607 : begin out <= 64'b1010100110100111101010101110001010011101000110101010100000010001; end
            14'd1608 : begin out <= 64'b1010100111001110101010011011011010101001100110110010100101111001; end
            14'd1609 : begin out <= 64'b1010100011010011001001001011011110100111000001001010001110001101; end
            14'd1610 : begin out <= 64'b1010011000101111101010101101100100100110011101010010101001110010; end
            14'd1611 : begin out <= 64'b1010010000100010100110011110010010100011001001000010101100001010; end
            14'd1612 : begin out <= 64'b1010011111001100101010000101100000101001011011101010011000101110; end
            14'd1613 : begin out <= 64'b0010011011111010101010100100101100011010110110000010100100101111; end
            14'd1614 : begin out <= 64'b0001111000110101101010011101111000011101110011100010011110001110; end
            14'd1615 : begin out <= 64'b0010101111101101101010001010111100101000110110011010100001011111; end
            14'd1616 : begin out <= 64'b0010010000111010001001110101000000101010011000001010101010101001; end
            14'd1617 : begin out <= 64'b1010100011011000001010110010111110101010110111101010100110000101; end
            14'd1618 : begin out <= 64'b0001111001111011001000010010100100100000010101100010010011100011; end
            14'd1619 : begin out <= 64'b0010101010111111101010001011100000101010111011000010101001000001; end
            14'd1620 : begin out <= 64'b0010010111010111101010100001001010101001001101101010101011111000; end
            14'd1621 : begin out <= 64'b1010011000001110101001001001100110101001110001010010100000010100; end
            14'd1622 : begin out <= 64'b1010100010000110001000111100100010010110111101100010011100110001; end
            14'd1623 : begin out <= 64'b1010100010010010001010100010100010100101000010001010100000011101; end
            14'd1624 : begin out <= 64'b1001110101111001101001110111100010101000011000010010100111011001; end
            14'd1625 : begin out <= 64'b0000011111001111001010001011001010100100101100110010011111011100; end
            14'd1626 : begin out <= 64'b0010100010110111101010000000001010101010101011101010100100100101; end
            14'd1627 : begin out <= 64'b0010101000000111100111110010110110100001000100111010010001000010; end
            14'd1628 : begin out <= 64'b0010100000111001101010100001000010100100001001111010001001100011; end
            14'd1629 : begin out <= 64'b1010101100011010001001110001110100101011110111100010101111100011; end
            14'd1630 : begin out <= 64'b0010101110111100101010100010010100011011100000101010100101001111; end
            14'd1631 : begin out <= 64'b0010011101101100001001001000000000100010010000011010001100111010; end
            14'd1632 : begin out <= 64'b0010101111101111001001111110010110100011101111011010101001100111; end
            14'd1633 : begin out <= 64'b1010010011110011001010110111010000100111111110011010100001011111; end
            14'd1634 : begin out <= 64'b1010100000110100100010101011110000100000000000101010101011011000; end
            14'd1635 : begin out <= 64'b0010001000011101101001011101111000100001111111001010011001011011; end
            14'd1636 : begin out <= 64'b1010101110011100001010110010110000101010111101100010010001000000; end
            14'd1637 : begin out <= 64'b1010100010101000001000010000010010101010111010101001111000011111; end
            14'd1638 : begin out <= 64'b1010101010100000101010110110010110101001101010000010101110101011; end
            14'd1639 : begin out <= 64'b0010000110000000001010111001000100100011111111101010101001101101; end
            14'd1640 : begin out <= 64'b1001110001101011101010000110000110100000101110101001111001100100; end
            14'd1641 : begin out <= 64'b1010011100001110100111101010011000101001010011011010101001011110; end
            14'd1642 : begin out <= 64'b1010101101011110001010100100110000101001010001000010100000110101; end
            14'd1643 : begin out <= 64'b1001110001000010001010101000111110011111110111111010100011101101; end
            14'd1644 : begin out <= 64'b1010100111010001001000101100000000100111110001001010101001000010; end
            14'd1645 : begin out <= 64'b1010001010000010001010011001111010101010100111001010100010001110; end
            14'd1646 : begin out <= 64'b0010010011000010000111001010001100101011101010100010000000110101; end
            14'd1647 : begin out <= 64'b1010100011110111101000111111011110100100111010001010010100101010; end
            14'd1648 : begin out <= 64'b1010011010001111100111000111100000011110111001011010011011010100; end
            14'd1649 : begin out <= 64'b1010000000101110101010011110100000101011101000101001000010111111; end
            14'd1650 : begin out <= 64'b1010100011010110001001000011010000101010100110000010100001111010; end
            14'd1651 : begin out <= 64'b0010101000100101001001000111010010100101111010000010011010001100; end
            14'd1652 : begin out <= 64'b0010101001000110101000110000111000100000101110101010011000110001; end
            14'd1653 : begin out <= 64'b0010011001111101001010111011110110101010110000000001101000011101; end
            14'd1654 : begin out <= 64'b0010101101101001101001000001111100101000110101001010010101010111; end
            14'd1655 : begin out <= 64'b0010001100000101001001011001111100101011111101101001111010110110; end
            14'd1656 : begin out <= 64'b0010100000101011001000110011111000101000000101111010101010101111; end
            14'd1657 : begin out <= 64'b0010100001110000001001111101010110100110000110110010101001111101; end
            14'd1658 : begin out <= 64'b1001111001100001101001101001000000101010101110010001111011001011; end
            14'd1659 : begin out <= 64'b1010101110010111100111100110100010100000000111101001111001011000; end
            14'd1660 : begin out <= 64'b1010100101110110001000110111100000011100111110100010101000101001; end
            14'd1661 : begin out <= 64'b1010100011010000000101111001101000100111101101100010101110111010; end
            14'd1662 : begin out <= 64'b0010101011001001001010011010101100100111101101100010100111010111; end
            14'd1663 : begin out <= 64'b0010010010011011001010000100001110101100000101000010010010001001; end
            14'd1664 : begin out <= 64'b1010001011110110001011000000000110100101000110000010101110110000; end
            14'd1665 : begin out <= 64'b0010100111111101001001101101000010101001100101000010100010110000; end
            14'd1666 : begin out <= 64'b1010101100001111000111101101100110100100001101101010001000100010; end
            14'd1667 : begin out <= 64'b1010010111010110100101011100000010100110110000101010100100011010; end
            14'd1668 : begin out <= 64'b0010101010101110001001010011000010100111100010101010011111111110; end
            14'd1669 : begin out <= 64'b0010010000101000101010110011110000100111111101011001000110111001; end
            14'd1670 : begin out <= 64'b1010100010110000001010001011101110101001001011000010001100100011; end
            14'd1671 : begin out <= 64'b1010100110011011001010101100100000011101010001001001101101110000; end
            14'd1672 : begin out <= 64'b1010101010001101001010010011001000101011010010111010100100001111; end
            14'd1673 : begin out <= 64'b1010011110011111100111111101100110100001010110000010001010110010; end
            14'd1674 : begin out <= 64'b1010100111011110101001011001010100100101000011111010100000101110; end
            14'd1675 : begin out <= 64'b1001111101100010001001101010001010101000100010110010010111110011; end
            14'd1676 : begin out <= 64'b1010100001111100001001110010101010011100100001101010100001101101; end
            14'd1677 : begin out <= 64'b1010011000001011001010111101101100101011100110100001111011110010; end
            14'd1678 : begin out <= 64'b1010101101010111100110000101011100100010000111110010100110011110; end
            14'd1679 : begin out <= 64'b0010101001001000001010111110011000101000100001011010010001010001; end
            14'd1680 : begin out <= 64'b0010101101101100100111101010110000011100111010011010010111101110; end
            14'd1681 : begin out <= 64'b0010100011001001000111011011010100101010001111111010101000011110; end
            14'd1682 : begin out <= 64'b0010101011101100001010010001101110100110001110000010101010000011; end
            14'd1683 : begin out <= 64'b0010100011100000001010100110000010011100110011101010100110110101; end
            14'd1684 : begin out <= 64'b1010101011100011001010111011111010100001001110011010101101011000; end
            14'd1685 : begin out <= 64'b0010100000101000001001100001111010101010010111111010010011001100; end
            14'd1686 : begin out <= 64'b1010101110011101001010010111110010101000100010101001101111011011; end
            14'd1687 : begin out <= 64'b1001100100110000101001110111011110100110010000101001110100011001; end
            14'd1688 : begin out <= 64'b1010101101100010101010101111110010100000100011111010010111100001; end
            14'd1689 : begin out <= 64'b0010010100000111101000101110110000100001100111010001100100011000; end
            14'd1690 : begin out <= 64'b1010100000011111101001011110101010100111000011111010010100110001; end
            14'd1691 : begin out <= 64'b0010000101010110101000010001111000101011101011110010011000100111; end
            14'd1692 : begin out <= 64'b0010100001000011101010000001011110100000001110111010101011001100; end
            14'd1693 : begin out <= 64'b0010101110000100001010100010101100100111010111011010011001101000; end
            14'd1694 : begin out <= 64'b0001110001110110000111010110011100101011111101110010011010010011; end
            14'd1695 : begin out <= 64'b0010100100001001101010111011010110100110001110101010001101111011; end
            14'd1696 : begin out <= 64'b0010010011001111101010101110100110101001101000011010101110000111; end
            14'd1697 : begin out <= 64'b0010011111101111000110101000110110101010100001011010010111001110; end
            14'd1698 : begin out <= 64'b0010000101110110101001111110001010101001110111001010011110001110; end
            14'd1699 : begin out <= 64'b1010100010100100101001111111010110101000111111000010100011111010; end
            14'd1700 : begin out <= 64'b1010100000110111001010101010010010100011001110111010010001101100; end
            14'd1701 : begin out <= 64'b1001110100110110001010100111000100011111010011110010001111101010; end
            14'd1702 : begin out <= 64'b0010000001110011101010010000000000010101111011101010001001011101; end
            14'd1703 : begin out <= 64'b0001111001100001101001110100110000100110000111111010100010000110; end
            14'd1704 : begin out <= 64'b0010100110011000001010110101010010100110111100101010001110000100; end
            14'd1705 : begin out <= 64'b1010100111011111001010011010100100101011010100100010011110111100; end
            14'd1706 : begin out <= 64'b1010101000010101001000110111010110100111011001111010001100010101; end
            14'd1707 : begin out <= 64'b1010101010100010001001111011101010100110000100111010010110111000; end
            14'd1708 : begin out <= 64'b0010101100010001001001110111111000101001100100111010000000110110; end
            14'd1709 : begin out <= 64'b1010101010110010001000001011001110100100001001010010101110111101; end
            14'd1710 : begin out <= 64'b0010100111010000101010110010100000101001001100101010101000110111; end
            14'd1711 : begin out <= 64'b0010100101001110101010101011011000101000000001110010001100011011; end
            14'd1712 : begin out <= 64'b1010101110001100001010101000000100101100001001011001110100100111; end
            14'd1713 : begin out <= 64'b1010011100110101100110011001110110100011110111100010010111111101; end
            14'd1714 : begin out <= 64'b0010101100001000101001011110000000100111001110110010110000001101; end
            14'd1715 : begin out <= 64'b1010100101100010101000010111101000101010100001110001111101101000; end
            14'd1716 : begin out <= 64'b0010100101110010001010110010101100100111100101100000010001100111; end
            14'd1717 : begin out <= 64'b1010101010000001001010010011100110101001001110000000100010001001; end
            14'd1718 : begin out <= 64'b0010101001000100101000110100100000100111010010101010000011001100; end
            14'd1719 : begin out <= 64'b0010101111100010001010000110101100101000010010111010100101011011; end
            14'd1720 : begin out <= 64'b0010100000100000001000110111110110101011110111100010101011101010; end
            14'd1721 : begin out <= 64'b0010011000111111001010011100111100101010010111110001101010001010; end
            14'd1722 : begin out <= 64'b0010010001000101001001001101010010011011101111010010101010111100; end
            14'd1723 : begin out <= 64'b0010101111000010101010100000011000101010110100010010000000101101; end
            14'd1724 : begin out <= 64'b0010000101100001101010010110010000100111001100101010000011000001; end
            14'd1725 : begin out <= 64'b1010101110101110101001100010100110101000110100111010001001011010; end
            14'd1726 : begin out <= 64'b0010101010001001001001010010111010101010101110000010001110111000; end
            14'd1727 : begin out <= 64'b0010101010110010001001001110001010100111001010001010000001111111; end
            14'd1728 : begin out <= 64'b0010010100000110100101001011010010100100100111001001111111100100; end
            14'd1729 : begin out <= 64'b0010100001100001101010010000001100011111110111000010000100000111; end
            14'd1730 : begin out <= 64'b0010100110101011101010101100011000100110001110100010101100101000; end
            14'd1731 : begin out <= 64'b0010101100010110100100000110110010101010010001001001110010010010; end
            14'd1732 : begin out <= 64'b1010011011101100101001110000110100101011111010011010100100100100; end
            14'd1733 : begin out <= 64'b0010101110111101001010100110111000100011111001011010101101010101; end
            14'd1734 : begin out <= 64'b1010010001001111001010110001100010100100110100111010010100010011; end
            14'd1735 : begin out <= 64'b1010100111100000001001111001001100101011110111111001100110111100; end
            14'd1736 : begin out <= 64'b1010101110010001101001011001100010101000000000110010101011111011; end
            14'd1737 : begin out <= 64'b0010100111010000101010110110000000100110001100011010101100010100; end
            14'd1738 : begin out <= 64'b0010100110000110001010100001010110101010000111101001110101001010; end
            14'd1739 : begin out <= 64'b0010010100100101001010100101110100100110010101010001011101011010; end
            14'd1740 : begin out <= 64'b0010011001110101100110001111000000101000100101001001101110100011; end
            14'd1741 : begin out <= 64'b1010010111001100101010000011110100101010101010100010000010000010; end
            14'd1742 : begin out <= 64'b1001101011010111101010110011000000101001010010000010000101100110; end
            14'd1743 : begin out <= 64'b1010011011110101101000001010001000101100000001111010011010011110; end
            14'd1744 : begin out <= 64'b1010100010000001001010010111111000100101111010011010100100111100; end
            14'd1745 : begin out <= 64'b0010100110010001001010110111100000011100110110001010100100111111; end
            14'd1746 : begin out <= 64'b1010000011001100101010110001000100101010001110100001110001101100; end
            14'd1747 : begin out <= 64'b0010100111000110001010111011100100011010001100100010101100100011; end
            14'd1748 : begin out <= 64'b0010011001010111101010011100011110101011111001001010010011001011; end
            14'd1749 : begin out <= 64'b0010011101001100101001100110001010100001011110011010000110101011; end
            14'd1750 : begin out <= 64'b1010011011110101001000000100010100100111100010111010101111101001; end
            14'd1751 : begin out <= 64'b1010101000001010101001111000111100100100000000101010010001011001; end
            14'd1752 : begin out <= 64'b0001100000100100101010111111011100101011111111011010011010100000; end
            14'd1753 : begin out <= 64'b1010101000101100001010100010011000101010010000111010101000110000; end
            14'd1754 : begin out <= 64'b0010011110101010001010100010100100101010011100010010100000010000; end
            14'd1755 : begin out <= 64'b1010101000111110001001010000111010100101010011010010101100101001; end
            14'd1756 : begin out <= 64'b0010100000100110101010011001000000101010000110010010101110100001; end
            14'd1757 : begin out <= 64'b1010011100010100101010010101001000010100111111111001100100001001; end
            14'd1758 : begin out <= 64'b0010001010011010001010001100011110100100010000111010000001110011; end
            14'd1759 : begin out <= 64'b1010101101100010101010110000001110010111100010101010101111011111; end
            14'd1760 : begin out <= 64'b0010100110000000101010011001101100101000100111001010011000000111; end
            14'd1761 : begin out <= 64'b0010101100101111001010110101011000100000001111011010011010111110; end
            14'd1762 : begin out <= 64'b1010011110101000101010010010011110101010011011011010100101001101; end
            14'd1763 : begin out <= 64'b0010100110010111101010111110001000101001110111000010101110000000; end
            14'd1764 : begin out <= 64'b1001100100010110001000101101110100100100101110111010011111110011; end
            14'd1765 : begin out <= 64'b0010011001000110000110001101101100101010000101111010100101100000; end
            14'd1766 : begin out <= 64'b0010101111111101001001110000011110101001011011111010100000100101; end
            14'd1767 : begin out <= 64'b0010100101001101001010100000000000100110101110110010001001010011; end
            14'd1768 : begin out <= 64'b1010011001000001101000001001110010101011101100111010100001010001; end
            14'd1769 : begin out <= 64'b1001010100011101101001100010011100011100011000011010100110101110; end
            14'd1770 : begin out <= 64'b0010100101100110000111000101110100100110110010000010100110000011; end
            14'd1771 : begin out <= 64'b1010010111101001101010001001011100101000001110100010010110010001; end
            14'd1772 : begin out <= 64'b1010100010010010101001111100111110100011000000110010011001001011; end
            14'd1773 : begin out <= 64'b1010100001101110001010100110110100001100000001011010011111100001; end
            14'd1774 : begin out <= 64'b1010100000111101101000001111000000011011010001011010100000001001; end
            14'd1775 : begin out <= 64'b0010001110110001001011000000000110100111111001101010000000111010; end
            14'd1776 : begin out <= 64'b0001011010001111101010001010101000000100001111011010011101100101; end
            14'd1777 : begin out <= 64'b0010011100111011001010100001011100100111010010101001111000001011; end
            14'd1778 : begin out <= 64'b0010100010111110101000000110100100010110011001011010101110011011; end
            14'd1779 : begin out <= 64'b0010100001100101000111011011001100011001111110111010101001000111; end
            14'd1780 : begin out <= 64'b1010100011011001000011111011100100100101110010100010101011001000; end
            14'd1781 : begin out <= 64'b0010010110101001001010111111010010100000111011011010100000100110; end
            14'd1782 : begin out <= 64'b1010101000111001101010110101110000100111011000110010100101111000; end
            14'd1783 : begin out <= 64'b1010100101100011100110101001100100101000000110011010101111110110; end
            14'd1784 : begin out <= 64'b0001101000011011101010011000000100001010011011000010100010001000; end
            14'd1785 : begin out <= 64'b1010010010011101001010010101011010101001110111111010100101011001; end
            14'd1786 : begin out <= 64'b0010011010000110101010000101111010101000010011000010100010000111; end
            14'd1787 : begin out <= 64'b1010010100001111001010010110010010011101001100010010011011011101; end
            14'd1788 : begin out <= 64'b1010101001011001101001100000100110101000010101000010010011000001; end
            14'd1789 : begin out <= 64'b0010011000111100101010110001000110100111111000101010010101000100; end
            14'd1790 : begin out <= 64'b1010101110101100001010010100001010100011001100010010101000111101; end
            14'd1791 : begin out <= 64'b1010100100110001001011000001101100100101001110000001110101000010; end
            14'd1792 : begin out <= 64'b1010101111101010001001111100101000101011001001101010101101110010; end
            14'd1793 : begin out <= 64'b1010101110111101101000011000100010100001010000111010001110100000; end
            14'd1794 : begin out <= 64'b0001100000001011101010001011011100101001011110010010101011001001; end
            14'd1795 : begin out <= 64'b1010100000010010000110011100110100100001001101100010101110001010; end
            14'd1796 : begin out <= 64'b1010100111000000001010011111101110101001010001011010101111010111; end
            14'd1797 : begin out <= 64'b1010101110100011100111111011000010101010100111111010100100001001; end
            14'd1798 : begin out <= 64'b1010101000100000101010010010101110100000100001110010100001011001; end
            14'd1799 : begin out <= 64'b0010101100101101001001011000110110101000001000111010011111111100; end
            14'd1800 : begin out <= 64'b0010010001100001001010111001111010101000010001001001111010100001; end
            14'd1801 : begin out <= 64'b1010001110110100001011000000101110101010011110110010100011101011; end
            14'd1802 : begin out <= 64'b1010100001101001101000101010000100101011101001101010101011110101; end
            14'd1803 : begin out <= 64'b1010101001000100100111000101000000101001100011001010010101011010; end
            14'd1804 : begin out <= 64'b0010101000000010101010011110101010101011000111101010011111101001; end
            14'd1805 : begin out <= 64'b0010010110001001101010001011011000100000001100100010100110111011; end
            14'd1806 : begin out <= 64'b0010100010100111101010100111100010100110011110110010001100010011; end
            14'd1807 : begin out <= 64'b1010100010111010001010011010000000101010000010001010000010100111; end
            14'd1808 : begin out <= 64'b1010101101110101101010010110101100010000001100010001110000000010; end
            14'd1809 : begin out <= 64'b1010101010000000000111010010010100101011010111000001110011110100; end
            14'd1810 : begin out <= 64'b0010001101101111101010110001001010100010101110001010100100111000; end
            14'd1811 : begin out <= 64'b1010001011000000101010101010001000100110000010111010100100110011; end
            14'd1812 : begin out <= 64'b1010101001010011000011100111010110011111001011001001111100110000; end
            14'd1813 : begin out <= 64'b0010100101011110001001100101101100100110110100110010000000111101; end
            14'd1814 : begin out <= 64'b0010101110011101001010110011000100101001001001011010101001101101; end
            14'd1815 : begin out <= 64'b0010100010111001001010000111100100101010110111010010100101001010; end
            14'd1816 : begin out <= 64'b1010011110100011101000010010110000011111111010000010011110011000; end
            14'd1817 : begin out <= 64'b1010001100010000001010011011101100101010110101001010100010010111; end
            14'd1818 : begin out <= 64'b0010100011111011101010111010001110101001100000001010100110101101; end
            14'd1819 : begin out <= 64'b0010011000000111001010111001011010101011011011101010100100000110; end
            14'd1820 : begin out <= 64'b1001111101010111101000111010011010101000111100101010100001000111; end
            14'd1821 : begin out <= 64'b0010100011000010101010110011101110100110100110101010100111011001; end
            14'd1822 : begin out <= 64'b0010101101010111101010011000010010101001010111110010100010100000; end
            14'd1823 : begin out <= 64'b1010010011100010101001000000101000101001010010100010011001011011; end
            14'd1824 : begin out <= 64'b0010010111111100101000000001100110101000000000011010011111000011; end
            14'd1825 : begin out <= 64'b1010011001110110101000000111011010100100010001101010011110100100; end
            14'd1826 : begin out <= 64'b0010100001010010101010101000011000101000100101110010101100111101; end
            14'd1827 : begin out <= 64'b1010010000011111001011000011111010101010010101111001011001000110; end
            14'd1828 : begin out <= 64'b1010000001000111001010110010101010101001101001100010100001110101; end
            14'd1829 : begin out <= 64'b0001111111100101001000011000000100100101001010011010101101010110; end
            14'd1830 : begin out <= 64'b0010100101000111000110101101100010100011011101101001010011100001; end
            14'd1831 : begin out <= 64'b0010001110010100101001101001011010101000110111100001110000011000; end
            14'd1832 : begin out <= 64'b1010011000001011001001101101100010100101001111010010100001010110; end
            14'd1833 : begin out <= 64'b0010101110100011101010000111001110100000010001101010001011000010; end
            14'd1834 : begin out <= 64'b1010100101101101101010010001011110010110101011111010010011001101; end
            14'd1835 : begin out <= 64'b1010100010111101001000000100111100100110100110101010101011101010; end
            14'd1836 : begin out <= 64'b1010100000111010000101011100001100101011001100111001110011100111; end
            14'd1837 : begin out <= 64'b1010100110100000001010001110010110101010010000110010100001000001; end
            14'd1838 : begin out <= 64'b1010010001010100001010110101011010011100100001100010011101000011; end
            14'd1839 : begin out <= 64'b0010100111010111001000000101001010100101110000001010011000000111; end
            14'd1840 : begin out <= 64'b1010100011110011101001010110000100101011001000010010001111000111; end
            14'd1841 : begin out <= 64'b0001111001011000101001010001011000101011001000000010100011011101; end
            14'd1842 : begin out <= 64'b1010101100111111101001000000011010100011000100011010100011001110; end
            14'd1843 : begin out <= 64'b1010101000011110001001001001011000100111000001100010101001101011; end
            14'd1844 : begin out <= 64'b1010101001011101001000101000100110101000110010100010100000000010; end
            14'd1845 : begin out <= 64'b1001110000111000101001111111110000100100011001000010100001001011; end
            14'd1846 : begin out <= 64'b0010010111111110101000100001101110101010010110100010010000011111; end
            14'd1847 : begin out <= 64'b1010101001100101000110011010000010100110110010110010011100110111; end
            14'd1848 : begin out <= 64'b1010100001100011001010110001000010010011110011110010010010000100; end
            14'd1849 : begin out <= 64'b1010011100001111000110010110010000100010001010000010101010010000; end
            14'd1850 : begin out <= 64'b0010010000101000001010011011101110100100001101000010101010011110; end
            14'd1851 : begin out <= 64'b0001111101110010001010000101000000101011001001101010101110100010; end
            14'd1852 : begin out <= 64'b0001111111000011101000110100111110101000011101011010010011011111; end
            14'd1853 : begin out <= 64'b0010000001100110000001111001011010101010001000111010101001110110; end
            14'd1854 : begin out <= 64'b0010101111000000101010110010100100101011111100000010000111010111; end
            14'd1855 : begin out <= 64'b1010101111100011001001110000011100100100001111011010010001111001; end
            14'd1856 : begin out <= 64'b0001011101011010001010111011100110100101010000100010100000110011; end
            14'd1857 : begin out <= 64'b0010100101011001001010001100010100100001001000100010010111001101; end
            14'd1858 : begin out <= 64'b1010010110101011001001101000011000100101000001010010101101011101; end
            14'd1859 : begin out <= 64'b1001010110010111101010101100010100101000001011000010100110011011; end
            14'd1860 : begin out <= 64'b0010101101001010001001101010010010100111110101000010011111100001; end
            14'd1861 : begin out <= 64'b1001110001110010001010011110100000100111011101110010011110101100; end
            14'd1862 : begin out <= 64'b1010011010110001001010101010001100101001101101110010010000010100; end
            14'd1863 : begin out <= 64'b1010000010111101001000111111111000101011000111100010011111001111; end
            14'd1864 : begin out <= 64'b1010100010011100000111111101111000101001101000001010101110100011; end
            14'd1865 : begin out <= 64'b1010100001000100001001111101110110101001101111011010100101000101; end
            14'd1866 : begin out <= 64'b1010101110001111101001011110101010100010101001111010011010010110; end
            14'd1867 : begin out <= 64'b0010010100110111101010000001001000011010100000101010010100010111; end
            14'd1868 : begin out <= 64'b1001110011000011101001100100000100101001010010010010001101010101; end
            14'd1869 : begin out <= 64'b1010010101010001101010011010011010101001100011010010011101000111; end
            14'd1870 : begin out <= 64'b0010101001110111101010010000001100100101010001111010011011010011; end
            14'd1871 : begin out <= 64'b0010100011101011001010110101100000100111001111111001000100010110; end
            14'd1872 : begin out <= 64'b1010101011111100001001111111010110101010101001101001110110011000; end
            14'd1873 : begin out <= 64'b0010000111011011101001111011000100100010001111010010001111101011; end
            14'd1874 : begin out <= 64'b0010100011011111001010100110011100100001011100011001110101110000; end
            14'd1875 : begin out <= 64'b1010011010110000001010100110011000101001000010101010110000110100; end
            14'd1876 : begin out <= 64'b1010011010101010101001100000000100100010101001001010010010011101; end
            14'd1877 : begin out <= 64'b1010100110101100101010100011111110101011111010111010101101000010; end
            14'd1878 : begin out <= 64'b0010100010011000001010101111110110101001010100010001100100110001; end
            14'd1879 : begin out <= 64'b1010011011111111101010110010011110100111010010100010101100010101; end
            14'd1880 : begin out <= 64'b1010100000011000001010011111001110101010101110011010100101011100; end
            14'd1881 : begin out <= 64'b1010100001001001101001001001011010101100000001111001000000000000; end
            14'd1882 : begin out <= 64'b0010100010011111101010101011100000100000110010000001111011000011; end
            14'd1883 : begin out <= 64'b0010000011100011100111101101010100101011000000100010100010001110; end
            14'd1884 : begin out <= 64'b0001111000000011001011000001000000100011110010111010000100101010; end
            14'd1885 : begin out <= 64'b1010000111110100001001011001011110101001010000100010101100011000; end
            14'd1886 : begin out <= 64'b0010100000111111101001100010011000101001011100011010001101000110; end
            14'd1887 : begin out <= 64'b1010101001011001101010100100111100100100010010010010001100000111; end
            14'd1888 : begin out <= 64'b1000111100011010101001101110111010101001011011001010101101101010; end
            14'd1889 : begin out <= 64'b0010100110101001001001011110001100100111101100010001100110000000; end
            14'd1890 : begin out <= 64'b1010011101000000001010101001101110101010000101101010100011010101; end
            14'd1891 : begin out <= 64'b0001111000111010001010111111000000101000111000101001111000110011; end
            14'd1892 : begin out <= 64'b0010000010100101101001001100100000011111110010111010101110011111; end
            14'd1893 : begin out <= 64'b1010100101000101001000100000110010101001111111010010100111101101; end
            14'd1894 : begin out <= 64'b0001110110111110001010100111111110100010001111101010100101111011; end
            14'd1895 : begin out <= 64'b0010000001110001101010111001000100011101100011101010011011001101; end
            14'd1896 : begin out <= 64'b0010101110110110101010110001001010100011100101000001110110100111; end
            14'd1897 : begin out <= 64'b1010101011010101101010001110101000100110111001100010100000110101; end
            14'd1898 : begin out <= 64'b0010100001011010001001011001101000101100000101100010101000101011; end
            14'd1899 : begin out <= 64'b1010010101001100101011000000011110101001101111100010011100010010; end
            14'd1900 : begin out <= 64'b0010011100110101101001011011111000100110110001001010101111100001; end
            14'd1901 : begin out <= 64'b0010010100110011001010101111010110100101111111010010100100011001; end
            14'd1902 : begin out <= 64'b0010001000101101101001010010001110101011111100010010101001010101; end
            14'd1903 : begin out <= 64'b1010100001111110101001101000001110100100100001100010001000111101; end
            14'd1904 : begin out <= 64'b1010010101001100001001100010001110101001101010000010000010011100; end
            14'd1905 : begin out <= 64'b0001101001011111001010111010110100101001100100000010001010010000; end
            14'd1906 : begin out <= 64'b1010010111110101101001011010011000101000011110001010100110010111; end
            14'd1907 : begin out <= 64'b0010010110110110001001010001011010100110111100011010100011001100; end
            14'd1908 : begin out <= 64'b1010011011101111101010111100011110101011111000111010101001101011; end
            14'd1909 : begin out <= 64'b0010011100111111100100110001110000101010001001101001110000011000; end
            14'd1910 : begin out <= 64'b1001110111111110001010100001101110101001101000000010100100001101; end
            14'd1911 : begin out <= 64'b1010101000101100001001010111111010101010000011000010010100100110; end
            14'd1912 : begin out <= 64'b0010100001000100101010001110011100101011101111001010100011110100; end
            14'd1913 : begin out <= 64'b0001000011011000101001011101011110101000100010111010101010101110; end
            14'd1914 : begin out <= 64'b0010010011000111101010000010001110100100111110011010101000001001; end
            14'd1915 : begin out <= 64'b0010100010011100001010011111100100100100100000100010010101111110; end
            14'd1916 : begin out <= 64'b0010101000111101101010101001010010011010111010111010100000010010; end
            14'd1917 : begin out <= 64'b1010100010100110100010001100111000011110110110110010011001000100; end
            14'd1918 : begin out <= 64'b0010010111010111001001110100011100101010001110001010100110100111; end
            14'd1919 : begin out <= 64'b1010000111100110101001001110011000101010100101001010001011111010; end
            14'd1920 : begin out <= 64'b1010010001111110001010011110010110101010110001001010101010011001; end
            14'd1921 : begin out <= 64'b1010101000001011001010000110111110011010000111100010100010101101; end
            14'd1922 : begin out <= 64'b1010011111000010001010000010010010100110001011010010010010000010; end
            14'd1923 : begin out <= 64'b0010011111011011001010110111011010100000111011000010100110100011; end
            14'd1924 : begin out <= 64'b1010100011000000100110110100011110101001000001100010101000000101; end
            14'd1925 : begin out <= 64'b1010100111010110001010100010111000011101000110100010100100000000; end
            14'd1926 : begin out <= 64'b0010011011111000001001100111011010011110100110110001111100110101; end
            14'd1927 : begin out <= 64'b0010101100111110000110000110010000101011000010001010110000111000; end
            14'd1928 : begin out <= 64'b0010100000001110001001001011100110100100000011111001000010100111; end
            14'd1929 : begin out <= 64'b0001011101111011101010100110100110100110011100010010011110001001; end
            14'd1930 : begin out <= 64'b1010101101011000001010111000111010100011011011000010011001011100; end
            14'd1931 : begin out <= 64'b1010010111100011001010100011001010101001111101011010011101101100; end
            14'd1932 : begin out <= 64'b1010010110110011001010001101111000101011000011001010101011110100; end
            14'd1933 : begin out <= 64'b0010101011010011101010100101000000011100000000011010011111000110; end
            14'd1934 : begin out <= 64'b1010011100110100101010000000110100101011010101011010100011110010; end
            14'd1935 : begin out <= 64'b1010010000101111001010110000001110011000011101000010011111101101; end
            14'd1936 : begin out <= 64'b1010100110011001101001000101100000101010010100111010000110110001; end
            14'd1937 : begin out <= 64'b0010010100010011101000000100011100100001001100010010000011110111; end
            14'd1938 : begin out <= 64'b1001111000011011101010100001101110100110100100011010000111111101; end
            14'd1939 : begin out <= 64'b0010001000001000101010100011011100101001000001110010100111111001; end
            14'd1940 : begin out <= 64'b0010010010110000001010101000111110100110100100101010100001000111; end
            14'd1941 : begin out <= 64'b1010011011101011000111111110011100101000111111000010010000001011; end
            14'd1942 : begin out <= 64'b1010011010010011101010001011111110101010000011001010100111010101; end
            14'd1943 : begin out <= 64'b0001100110001111101000101011001010100110011011101010011100011110; end
            14'd1944 : begin out <= 64'b0010101011001100001010100011001010101010110001010010001011001011; end
            14'd1945 : begin out <= 64'b1010001010101100001010100001111010101000001001101010100001110011; end
            14'd1946 : begin out <= 64'b0010100001110110001010001010011010100000101110100010100111001001; end
            14'd1947 : begin out <= 64'b1001110000001101001001111000101000101001000010100010100111101011; end
            14'd1948 : begin out <= 64'b1010100010101001101001001110100010101001110011110010011011111110; end
            14'd1949 : begin out <= 64'b0010011000010110100100111011011100100100110100111010101011110111; end
            14'd1950 : begin out <= 64'b0010101011010100001010110000101100101010010011100010110001001011; end
            14'd1951 : begin out <= 64'b0010010110010001101010010011101000101010010010101010010111011111; end
            14'd1952 : begin out <= 64'b0010000010111001100011001010101110101010111101110010101100000101; end
            14'd1953 : begin out <= 64'b1010100110001000001010110110010000100110011111001010010111100011; end
            14'd1954 : begin out <= 64'b1010011111110011001010110111111100100011000000011010101100010010; end
            14'd1955 : begin out <= 64'b1010011110110001000110101101111110100101101100000010011100000101; end
            14'd1956 : begin out <= 64'b0010101100001110101010010011100100010101011000101010001111101010; end
            14'd1957 : begin out <= 64'b1010101010100101101001000001010000101010000011001010010001101001; end
            14'd1958 : begin out <= 64'b1001101111001010100111100011010000101011101001001001100110111010; end
            14'd1959 : begin out <= 64'b1010000110010111001010001110001110101001111001110010001101011010; end
            14'd1960 : begin out <= 64'b1010100011001001101010011101101110101001001011011010000010010011; end
            14'd1961 : begin out <= 64'b0010100100000100101000000011100110100001001000001010100011011010; end
            14'd1962 : begin out <= 64'b1010100100001000101010110100101100101000011101000010100110111100; end
            14'd1963 : begin out <= 64'b1010100111110110101010100111100100011010100110100010010110110100; end
            14'd1964 : begin out <= 64'b0010011011111011001010111001100110100111000111101010000110110011; end
            14'd1965 : begin out <= 64'b0010101000111011101010101111010110011111000111011010010000010011; end
            14'd1966 : begin out <= 64'b1010101011001111100111100011101100101000111011100010110000100001; end
            14'd1967 : begin out <= 64'b0010100101011011101010110110011100100010111111111010101101001001; end
            14'd1968 : begin out <= 64'b0010010011111110101010010111011110100010100010100010100010101100; end
            14'd1969 : begin out <= 64'b0010011100001010101010011100001010011110100101000010000111011011; end
            14'd1970 : begin out <= 64'b1001110011011100101001111110010000101000101001000010101101111110; end
            14'd1971 : begin out <= 64'b0010101001111011101010101010011100100100101010010010100011100001; end
            14'd1972 : begin out <= 64'b0010100000001000001010101100010100100011000011011010101000100010; end
            14'd1973 : begin out <= 64'b1010101000101111101010101000010110100001100110100010100001011011; end
            14'd1974 : begin out <= 64'b0010011111010110101001000110010100100101010010010001000011000100; end
            14'd1975 : begin out <= 64'b1010100010001101001010100001100010100111000111000010011100101100; end
            14'd1976 : begin out <= 64'b0010011010011010101010000000101000100100010010011010110001101100; end
            14'd1977 : begin out <= 64'b1010100001111001001010010100000000100100000000101010011001100000; end
            14'd1978 : begin out <= 64'b1010001001110011101010010110011100101001001100001001111010010101; end
            14'd1979 : begin out <= 64'b1010101001011100101010100100011110101000011110000010100000010010; end
            14'd1980 : begin out <= 64'b0010010100101110101010100001100110101010011101111000110101011110; end
            14'd1981 : begin out <= 64'b0010101100111111001001101011001100101001000111010010100000011000; end
            14'd1982 : begin out <= 64'b0010000001011111001001001101111000001110011010010010101101010100; end
            14'd1983 : begin out <= 64'b1010100101011000101000111001010000101011001110011010010101001101; end
            14'd1984 : begin out <= 64'b0001101011001100001010100001000110100010110100101010010111001111; end
            14'd1985 : begin out <= 64'b1010000010100101000111010101111010100010110110011010001011001111; end
            14'd1986 : begin out <= 64'b1010101011100101101001100001100110101011000100110010101101111011; end
            14'd1987 : begin out <= 64'b0010100011111100001001100111101010101000011001010010010000101101; end
            14'd1988 : begin out <= 64'b1010011010010100001000010110000010100111010011110000110111000001; end
            14'd1989 : begin out <= 64'b1010100111010100001010010100110110101000000101110010100100011101; end
            14'd1990 : begin out <= 64'b1010100110100110001001101101100100101010110010111010100000000011; end
            14'd1991 : begin out <= 64'b0010010111111011101010001110111110101001101100110010010010001111; end
            14'd1992 : begin out <= 64'b1010100100100001101010001000010110101011000111000010100111100100; end
            14'd1993 : begin out <= 64'b1001110100100001001001111010111110100101101100101010100001111001; end
            14'd1994 : begin out <= 64'b0010000000000001001010101101101110011000000011001010010001011101; end
            14'd1995 : begin out <= 64'b0001111000011100101001001000000110101010000010010010101010110101; end
            14'd1996 : begin out <= 64'b0010100111001010100111100101100010100111100001101010010100001000; end
            14'd1997 : begin out <= 64'b0001100010001010101000101011011010101000011111100010011101010111; end
            14'd1998 : begin out <= 64'b1010101101010001101001011001010000101010011101111010010100110101; end
            14'd1999 : begin out <= 64'b0010000111011011101010101111000100101001101010000010100110010111; end
            14'd2000 : begin out <= 64'b0010100001001110001010000101001110100011111011011010000011101100; end
            14'd2001 : begin out <= 64'b1010101010011011001000010000001010101010000011000010011011010101; end
            14'd2002 : begin out <= 64'b0010101100101100101001111001001000100001011000111010011110101001; end
            14'd2003 : begin out <= 64'b0010100101000000100111100101010100101001010101010010101100100101; end
            14'd2004 : begin out <= 64'b0010101100101110101000010100000010101010111001000010101001010011; end
            14'd2005 : begin out <= 64'b0010100010100111101010001011111000101010001010101010100011010000; end
            14'd2006 : begin out <= 64'b1010011000111111001010110001011010100001000010001010100110010010; end
            14'd2007 : begin out <= 64'b1010001100010110100111000100100110101000000111010010001011001010; end
            14'd2008 : begin out <= 64'b0010101111101110001010110101001000010101110000100010010011000000; end
            14'd2009 : begin out <= 64'b0010100010111001001010101101000000011000111000001010011001001101; end
            14'd2010 : begin out <= 64'b1010001001000010101010001000000000100100111111100010100110100010; end
            14'd2011 : begin out <= 64'b1010010110111111001010000111101000100000110011100010011100011110; end
            14'd2012 : begin out <= 64'b0010001011010101101001110100010010001111110011100001110000100010; end
            14'd2013 : begin out <= 64'b1010100101100011001010110101110000101000001101001010100111001100; end
            14'd2014 : begin out <= 64'b0010100000010010000111011100011100100101000000100010000101001100; end
            14'd2015 : begin out <= 64'b0010100001100100001010010100010110100110011000101010101000011101; end
            14'd2016 : begin out <= 64'b1010011100010010100110010111100010011101001100101010010011101000; end
            14'd2017 : begin out <= 64'b1010010100000111001010101110111010101000101011100010001000101110; end
            14'd2018 : begin out <= 64'b1010101101101100101001010010101010100100000110001010101100101101; end
            14'd2019 : begin out <= 64'b0010010101100111001010001111001010101001101110011010100100011111; end
            14'd2020 : begin out <= 64'b0010010111111011001001110111110100010110100100011010101010000001; end
            14'd2021 : begin out <= 64'b1010011011011000000111101011100100100000001000001010100000001110; end
            14'd2022 : begin out <= 64'b1010101101011101001010001100010100101000011000010001110011111010; end
            14'd2023 : begin out <= 64'b0010101110101000001010110000101000100000011111000010101011110101; end
            14'd2024 : begin out <= 64'b0010000000100010100101110001000010101010101111010010001000101111; end
            14'd2025 : begin out <= 64'b1010101011001011101001110001110100101001011100100010100001011101; end
            14'd2026 : begin out <= 64'b0010100100111111101001110110010000101001100010010010100000100000; end
            14'd2027 : begin out <= 64'b1010010101111111101001000110111010100110110100110010011110111010; end
            14'd2028 : begin out <= 64'b1010010001011100001011000001100110100101011101110010100110100001; end
            14'd2029 : begin out <= 64'b0010010100010110101010000100001010101011110011010010100001111000; end
            14'd2030 : begin out <= 64'b1010100011011110101010101111011010100111010001000010101001110001; end
            14'd2031 : begin out <= 64'b0010010100001011101000111010011000101011100001101010100011001101; end
            14'd2032 : begin out <= 64'b1010100111111110101010101000111010011100010011000010011111001000; end
            14'd2033 : begin out <= 64'b0010100101011110001010100100110110101001110110010010100100010011; end
            14'd2034 : begin out <= 64'b0010100001110100001010001001000010011110110000100010100101001111; end
            14'd2035 : begin out <= 64'b1010101111001111101010011101111010100101011011011010010001111000; end
            14'd2036 : begin out <= 64'b1010000101011011001010000000000000101000000011110001111011111110; end
            14'd2037 : begin out <= 64'b0010100000111110001010011010010000100010101010100010010100000011; end
            14'd2038 : begin out <= 64'b1010000111101111000111010001011100010000111010001010011011001000; end
            14'd2039 : begin out <= 64'b1010101000111011001000010001000010101010110001111010100111110101; end
            14'd2040 : begin out <= 64'b0010000111101011101010001101001010101011110111101010101111000101; end
            14'd2041 : begin out <= 64'b1010100001110101101010111011010100011101110111100010101110110001; end
            14'd2042 : begin out <= 64'b0010100010110110001010110001100110101010000001010010010000101000; end
            14'd2043 : begin out <= 64'b1010100110001000101001101101000000101001101111000010100101100111; end
            14'd2044 : begin out <= 64'b1010100100001010001001001011000010011010010100011010000110101110; end
            14'd2045 : begin out <= 64'b1010100111011101101001100111111000100101100001101010100010010111; end
            14'd2046 : begin out <= 64'b0010100001001010001000010110011010100011011001000010100110100100; end
            14'd2047 : begin out <= 64'b1010101001110100001000001000011110101010100111000010100111000101; end
            14'd2048 : begin out <= 64'b1010101101000111001010000111100100101001000111100010000000001110; end
            14'd2049 : begin out <= 64'b0010100101110111001000001110001110101001100000111010100001101010; end
            14'd2050 : begin out <= 64'b1010011011110100001010011010001000100000100110011010100000111100; end
            14'd2051 : begin out <= 64'b1010101011111100101010011011010110011000011101000010101010111111; end
            14'd2052 : begin out <= 64'b1001100011001110101010111000011000100010110000011010011101110001; end
            14'd2053 : begin out <= 64'b0010100001001110001000011001100110101011110010111010001100110011; end
            14'd2054 : begin out <= 64'b0010011010001011101010100110010110100101001100011010001010000101; end
            14'd2055 : begin out <= 64'b0010100110010010001010101110001000101001101111011010101110101010; end
            14'd2056 : begin out <= 64'b0001110101011100001010110101100100101000111001110010101001001011; end
            14'd2057 : begin out <= 64'b0010001010100110101010111010001110101001101100001010010111010111; end
            14'd2058 : begin out <= 64'b0010101101011010001010011010011000011011010101001010100110000111; end
            14'd2059 : begin out <= 64'b1001110100100001101010011010110100101000111111100001000011001010; end
            14'd2060 : begin out <= 64'b0010100101110000001010001111010100100010100110100010101101100000; end
            14'd2061 : begin out <= 64'b1010101100110011001010110110010110101001111100111010000010010010; end
            14'd2062 : begin out <= 64'b0010011101001111001010011100001110100001001011011010101111001010; end
            14'd2063 : begin out <= 64'b0010100101110100001001000111101100100100011001110001111100101100; end
            14'd2064 : begin out <= 64'b1010100110100111001010010011110110100011000010000010101000010101; end
            14'd2065 : begin out <= 64'b0010000100010100001010101011000000100101110000011010100001101111; end
            14'd2066 : begin out <= 64'b0010100001101011101000011110010000101001111111011010100010010101; end
            14'd2067 : begin out <= 64'b1001110110100110101010111010110000101011101110011010101101001100; end
            14'd2068 : begin out <= 64'b1010100001010110001010110000100000011111010110011010100010000001; end
            14'd2069 : begin out <= 64'b1010100101001101101010110111100000101001110111000000000001111110; end
            14'd2070 : begin out <= 64'b1010101011111111001001110011001000101010001111111010010111011100; end
            14'd2071 : begin out <= 64'b0001110111110011101010000001010000101010011011011010011101101111; end
            14'd2072 : begin out <= 64'b0001011111000101001001001101011010011111001111110010100100000011; end
            14'd2073 : begin out <= 64'b1010010110001101101010000011110000101011110010111010101001010010; end
            14'd2074 : begin out <= 64'b1010101101110011001001011000110100101010010001100010010100101100; end
            14'd2075 : begin out <= 64'b0010101000110101001010011110100010101010110101010010011101100101; end
            14'd2076 : begin out <= 64'b1010000011101111001010001101101000100100100111110010101000101111; end
            14'd2077 : begin out <= 64'b0010000110000100101010101100110110100000111110100010101010000001; end
            14'd2078 : begin out <= 64'b1010011100110001001000100111000000100110010001110010100101011100; end
            14'd2079 : begin out <= 64'b1010100101101100101010110011010100011001000100011010000011001111; end
            14'd2080 : begin out <= 64'b0010011001101110101010001101100110100101000100101010010011010111; end
            14'd2081 : begin out <= 64'b1010100001010100001010111100011110011111111001000010100101110011; end
            14'd2082 : begin out <= 64'b1010101001001111101010111001010100101000101001111010100011010011; end
            14'd2083 : begin out <= 64'b1010100011001101101010010101001110101001111111101010100011010001; end
            14'd2084 : begin out <= 64'b1010010010110111001001011000000000101011001100101010000001000001; end
            14'd2085 : begin out <= 64'b0010101010101100100111101110000110101011011111101010001101100011; end
            14'd2086 : begin out <= 64'b1001111000111110001001111001000010101010001010000010100111010101; end
            14'd2087 : begin out <= 64'b1001110001100010001001000101110110101011000110111010101001100011; end
            14'd2088 : begin out <= 64'b1010101100101011001010100010110100101010101101000010000110001010; end
            14'd2089 : begin out <= 64'b0001110110100100101001100000000110101011010111011010000110111010; end
            14'd2090 : begin out <= 64'b0010011001100011001010110101010110011110100001111001101010111100; end
            14'd2091 : begin out <= 64'b1010100100111100101000110000000000101010100000100010010101001100; end
            14'd2092 : begin out <= 64'b1010010110101000101001000011000000100111100000011010100101111001; end
            14'd2093 : begin out <= 64'b0010101101010001001001000100111100101011001110110010011111101100; end
            14'd2094 : begin out <= 64'b0010000000110111000111101111111100101001100111111010010010001110; end
            14'd2095 : begin out <= 64'b0010100100110010101001001011000010101011101001111010001010100110; end
            14'd2096 : begin out <= 64'b1010101100111111101010000111110000101001100100010010101011101011; end
            14'd2097 : begin out <= 64'b1010010100110111101010011110111010100101000010110010011000100001; end
            14'd2098 : begin out <= 64'b1010100100011101001010110001001110010101111011000010000111010111; end
            14'd2099 : begin out <= 64'b0010011011101111100110100010000010100101011011000010100011100010; end
            14'd2100 : begin out <= 64'b1010101011111010001001101111000100101010111011100010010100010001; end
            14'd2101 : begin out <= 64'b1010011001011111001010100111001010010110101110110010100101000001; end
            14'd2102 : begin out <= 64'b0010010001000000101001011011000110100100000111011010100010001010; end
            14'd2103 : begin out <= 64'b1010010001001111101010111110010100101001110010101001111010011011; end
            14'd2104 : begin out <= 64'b1001110111110001100111000010100110100110001011011010100001010101; end
            14'd2105 : begin out <= 64'b1010011011101110101010001001011110101010110010101010101110101110; end
            14'd2106 : begin out <= 64'b1010010011111000101010000010100100101010111001101010101110111011; end
            14'd2107 : begin out <= 64'b1010001001110011101010101110010110101000101010101010010100111010; end
            14'd2108 : begin out <= 64'b0010100100111101001010101011101110101011110110010010000101111010; end
            14'd2109 : begin out <= 64'b1010101110111110101010010101000000101000011100010010100110010010; end
            14'd2110 : begin out <= 64'b1001111001011000001010010110110010011010111111011001110011111010; end
            14'd2111 : begin out <= 64'b1010100000110010100111011000001010011011011010011010100000110101; end
            14'd2112 : begin out <= 64'b0001000000010011001001100100100000100111100001101010001011000000; end
            14'd2113 : begin out <= 64'b1010001100010010101001101110101110101000000010110010100001010001; end
            14'd2114 : begin out <= 64'b1010100000100110001010011000010010101011110001101010001110110100; end
            14'd2115 : begin out <= 64'b1010100111100111001000001111000110101000110100111010101000001001; end
            14'd2116 : begin out <= 64'b0010100000111110001001000001111100001100011100000010101110101011; end
            14'd2117 : begin out <= 64'b0010010100000010000111110001101010101000110011100010001100100101; end
            14'd2118 : begin out <= 64'b0010101011001101101010110010000000101000110011110010101111000101; end
            14'd2119 : begin out <= 64'b1001110111111110101001011110111000101001000001001001110101101111; end
            14'd2120 : begin out <= 64'b0010010100001010000101101111000010101001101010101010100101110100; end
            14'd2121 : begin out <= 64'b0010101110110101101001110101111000100110110011011010010110101011; end
            14'd2122 : begin out <= 64'b1010101010110000001001100111010110100101011001101010011000100000; end
            14'd2123 : begin out <= 64'b1010010011101101001000011110001110101001011011111010101110100101; end
            14'd2124 : begin out <= 64'b0010100001100101101010011011100100011100011000111010101010111001; end
            14'd2125 : begin out <= 64'b0010100100101111001001001011000010100100001011000010010011111110; end
            14'd2126 : begin out <= 64'b0010101100010000100111111110001100101001000010001010010010100001; end
            14'd2127 : begin out <= 64'b0010101110000110001001100011110010100110011110110010010001000010; end
            14'd2128 : begin out <= 64'b0010001111011110001010101000010000100110000011111001111000110100; end
            14'd2129 : begin out <= 64'b1010100101001100101001000100101100100100001100011010100001100011; end
            14'd2130 : begin out <= 64'b1010100001000011000111010110100100101011010110100010101111110010; end
            14'd2131 : begin out <= 64'b0010100100110011001010110101001010101001000111111001101010111011; end
            14'd2132 : begin out <= 64'b1010011111001100001010001001000010100001100010000010000010100010; end
            14'd2133 : begin out <= 64'b0010101111000111100110011111001000101011100100100001100100000111; end
            14'd2134 : begin out <= 64'b1001111101000001101010111101111110100011011001101010000000001100; end
            14'd2135 : begin out <= 64'b0010101001100010101001000100100000101001111110100010001001100110; end
            14'd2136 : begin out <= 64'b0001110010100111101001111111111100011001001110010010101011100110; end
            14'd2137 : begin out <= 64'b1010101010110011001001110100011110100110111010100010101110111010; end
            14'd2138 : begin out <= 64'b0010010011001100001010001101111000100110000010100010000011010011; end
            14'd2139 : begin out <= 64'b0010101110100010101001011101110110100101011011011010011100100110; end
            14'd2140 : begin out <= 64'b0010010100100010001001001111011100101011001111001010010001110110; end
            14'd2141 : begin out <= 64'b1010101001110111001010100101010010100000110010010010011001101111; end
            14'd2142 : begin out <= 64'b0010011110011110001010110001100110100110111001100010010100110110; end
            14'd2143 : begin out <= 64'b0010100001101111100100010110001100101011011011011010100101111100; end
            14'd2144 : begin out <= 64'b1001100011001001101010000011101110100010100000001010100000011111; end
            14'd2145 : begin out <= 64'b1010000001010000100111111101101100101001010010101010011101001011; end
            14'd2146 : begin out <= 64'b0001110010101011001000101111101100100100010010010010001110111101; end
            14'd2147 : begin out <= 64'b0010000101010001100101100100100000101000111110100001110011011101; end
            14'd2148 : begin out <= 64'b0010010100010000101010110100000110101001010110001010010111101110; end
            14'd2149 : begin out <= 64'b1010101100011111101010101111000110100000010001101010101100110010; end
            14'd2150 : begin out <= 64'b1010101111100110001010110001100010101011110111001010100010000110; end
            14'd2151 : begin out <= 64'b0001111101000110001010010011100000101010100100111010011001010001; end
            14'd2152 : begin out <= 64'b0010100101011111001010000110111000101000011100111010101111000111; end
            14'd2153 : begin out <= 64'b0010011101100001001000001001011000101011010110011010100101110101; end
            14'd2154 : begin out <= 64'b1010100011000001001010110110001000101011110100110010100100101100; end
            14'd2155 : begin out <= 64'b0010011101010011001001100111100110100101001001000010101110111000; end
            14'd2156 : begin out <= 64'b0010000010101011000110110001011010100010010001010010000111100110; end
            14'd2157 : begin out <= 64'b0010100110001011000111000111101010101010100001110010100010101010; end
            14'd2158 : begin out <= 64'b0010100110111010001010000000010110101011001101111001010100000001; end
            14'd2159 : begin out <= 64'b1010100000100000001001101101110010100111110110101010100001110100; end
            14'd2160 : begin out <= 64'b1010100000110000001001001101010110100111010101111010101011101110; end
            14'd2161 : begin out <= 64'b1010100011000011101010001001010010100101100110101010100001101001; end
            14'd2162 : begin out <= 64'b1010011000011110101010101001101010011110000011110010011001010111; end
            14'd2163 : begin out <= 64'b1010100101000100001010000110101010100100101110101010100011000101; end
            14'd2164 : begin out <= 64'b1010101011100100101010011110000100100101111100101010011010001111; end
            14'd2165 : begin out <= 64'b1010100111000010001000000011001000101011101101011010100100010101; end
            14'd2166 : begin out <= 64'b0010010000011111001010111011000100100110100001010010100110011111; end
            14'd2167 : begin out <= 64'b0010101001100101101010001100101110100101101101111010101011001000; end
            14'd2168 : begin out <= 64'b0010010001101110001010011111100100100101110011100010101100001110; end
            14'd2169 : begin out <= 64'b1010101001111001001001110001101000100101111011011010011010011101; end
            14'd2170 : begin out <= 64'b1010010001111010100111011000111010101011111000111010100001100010; end
            14'd2171 : begin out <= 64'b0010001111010111001010001101010100101011011000000001111000101100; end
            14'd2172 : begin out <= 64'b1010100000111100100110101011101100100110100101000010010011011110; end
            14'd2173 : begin out <= 64'b0010100101101001001001000000100000100100001001010010101111001000; end
            14'd2174 : begin out <= 64'b1010100011010110001010001000110010100101010101100010100001101101; end
            14'd2175 : begin out <= 64'b1010101101101001100111011000000100100111101100000010011001001101; end
            14'd2176 : begin out <= 64'b0010011111110011001010101100011000101000100110000010101110010110; end
            14'd2177 : begin out <= 64'b0010100111110101101010101000011010101010101101010010100000001110; end
            14'd2178 : begin out <= 64'b0010100001110100100111000111111010011100000100010010100101001010; end
            14'd2179 : begin out <= 64'b0010010001110100001010101111000000101010111000110010101111100010; end
            14'd2180 : begin out <= 64'b1010101101100100101001000010011110100001110000011010001111101100; end
            14'd2181 : begin out <= 64'b1010000101000010001010101110110010100110001011111010001000100101; end
            14'd2182 : begin out <= 64'b1010001000001100001001010000111000100111101100011010100100100101; end
            14'd2183 : begin out <= 64'b1010011001000000001010110101001100100111011011010001100100100110; end
            14'd2184 : begin out <= 64'b1001101000010011101001111010000110011100010010010010011001101001; end
            14'd2185 : begin out <= 64'b0010100001001010101010101010101000100111010100101010101011110001; end
            14'd2186 : begin out <= 64'b0010001001001110101010101010111010101001010011010010101111000011; end
            14'd2187 : begin out <= 64'b0010010011011111101001110000110110101011110100101010100001111100; end
            14'd2188 : begin out <= 64'b0010101110000111101010111111100010100111110011111010010011010010; end
            14'd2189 : begin out <= 64'b0010101110101100001010010011101100100010000110000010100010010111; end
            14'd2190 : begin out <= 64'b0010000001111111001001111000010010101001001001110010101110001010; end
            14'd2191 : begin out <= 64'b0010010010101010001001001110000000011010111001100010101110010110; end
            14'd2192 : begin out <= 64'b0010101011110111001010110010101010100001111100101010101000111100; end
            14'd2193 : begin out <= 64'b1001100101010010100101101011101110100110011001111010100100010010; end
            14'd2194 : begin out <= 64'b0001111010001010101010011001110010101011110100100010100100111000; end
            14'd2195 : begin out <= 64'b1000100010001001001000111111011010100100110111111010010100100101; end
            14'd2196 : begin out <= 64'b1010100110011111001010100000100000100100100111010001101011000000; end
            14'd2197 : begin out <= 64'b1010101100101110101001001010100110101011100000101010001000011000; end
            14'd2198 : begin out <= 64'b0010100111110001101010001011100010100100110111001010101001000000; end
            14'd2199 : begin out <= 64'b0010101100100101001010110110001010101010000001000010010100100110; end
            14'd2200 : begin out <= 64'b1010100011001001001000100100011000101001100101010010100000010011; end
            14'd2201 : begin out <= 64'b0001010100010110101010100110011010101011111010100010100100100101; end
            14'd2202 : begin out <= 64'b1001100000010111001001110011011000101011110100101010100000100100; end
            14'd2203 : begin out <= 64'b0010100111001011101000010111111010100001111101100010010011100111; end
            14'd2204 : begin out <= 64'b1001100010110111001010111000011110011001010011110010100010000111; end
            14'd2205 : begin out <= 64'b1010100000100010000111110010010100101001010001101010010001000101; end
            14'd2206 : begin out <= 64'b0010100011101100001010100100101100100101110001011010100010110010; end
            14'd2207 : begin out <= 64'b1001101000111000101000111001000000100100110001110010001111110100; end
            14'd2208 : begin out <= 64'b0010101010100100001001010011001110100110000101011010101010000111; end
            14'd2209 : begin out <= 64'b0010010110010100001000101011101010101011000010110010000010001011; end
            14'd2210 : begin out <= 64'b0010001101011110001001001010101110100100010000000010010100011010; end
            14'd2211 : begin out <= 64'b0010001111011000001001101101001110100010011000001010010100101000; end
            14'd2212 : begin out <= 64'b1001110011110000001010010010101000100111011000001010011000000111; end
            14'd2213 : begin out <= 64'b1010100101001110000111001010011010101001101001011010101011101010; end
            14'd2214 : begin out <= 64'b0010101100001110101010110111110110100111101011011010011110110101; end
            14'd2215 : begin out <= 64'b0010010101110110101010100000101000100011010011011010101100111000; end
            14'd2216 : begin out <= 64'b1010010100000001101010100010101110101001000000001010001111011000; end
            14'd2217 : begin out <= 64'b1010010100001111001010000010101000101010011110111010100110011000; end
            14'd2218 : begin out <= 64'b0010101110010110001010110100101010101010110000110010101010100111; end
            14'd2219 : begin out <= 64'b0010010100100110101001111010100010011000001111011010101010011110; end
            14'd2220 : begin out <= 64'b0010100011101100001001101011000110100111001110011010100000001011; end
            14'd2221 : begin out <= 64'b0010000000100010000101110110101100101010101011110010001101011110; end
            14'd2222 : begin out <= 64'b1010101001110001101010000100000100100110010000001010100011000011; end
            14'd2223 : begin out <= 64'b1010001010111011101010100111000110100101010001100010000111100101; end
            14'd2224 : begin out <= 64'b0001110010101000101001110100001010100011111100001010100011000000; end
            14'd2225 : begin out <= 64'b0010101100001100101001111001101000100100011001111010011001101101; end
            14'd2226 : begin out <= 64'b0010100111011011101001110111001010100001000010100010001000110011; end
            14'd2227 : begin out <= 64'b0010101110100101001010101100101010100100000101111010101001101110; end
            14'd2228 : begin out <= 64'b0010101110110101100101001010000100100100010101101010000000010001; end
            14'd2229 : begin out <= 64'b0010011010001100100101010110001000101011000011110010101010100101; end
            14'd2230 : begin out <= 64'b0010101101101010001010111001000000100111010001011010101011000100; end
            14'd2231 : begin out <= 64'b0001111101010101101000111101000110101010000111001010010101101100; end
            14'd2232 : begin out <= 64'b1010011000000111001010000101011110101010001111100010011110111010; end
            14'd2233 : begin out <= 64'b1010100100100011001010011011001000101010011110101010100101110000; end
            14'd2234 : begin out <= 64'b0010011101011001101000111111100110101001101110111010100001110010; end
            14'd2235 : begin out <= 64'b1010101010011101001010001011001000100111011101111010000000000000; end
            14'd2236 : begin out <= 64'b1010101100100010101010101100001000101010010000110010010101000101; end
            14'd2237 : begin out <= 64'b1010101100011000101010010001100100100100111110110010010110111011; end
            14'd2238 : begin out <= 64'b0010011000010001100111001001100110101001111101000001100000011111; end
            14'd2239 : begin out <= 64'b0001111000100100101001001011100100100001011000101010101110111101; end
            14'd2240 : begin out <= 64'b0010101010110101101010101011111000101011001011110010100111100001; end
            14'd2241 : begin out <= 64'b0010100111110110001010010000110000101000010100010010100101110001; end
            14'd2242 : begin out <= 64'b1001111111000101100101010100000010101011111110011001111101011110; end
            14'd2243 : begin out <= 64'b0001111100110110101010110101000100010101000000101010100001011110; end
            14'd2244 : begin out <= 64'b0010101001001111101010011100011110100010010110101010100101111100; end
            14'd2245 : begin out <= 64'b0010010001111001101000110111101000101001110001010010010111100001; end
            14'd2246 : begin out <= 64'b1001100000011011101000111000111010100101100000110010100110111100; end
            14'd2247 : begin out <= 64'b1010010100100111101000111110010110100100010011000010010110111011; end
            14'd2248 : begin out <= 64'b0010101010110001100111011100101100101011011010100010101001110111; end
            14'd2249 : begin out <= 64'b1010000111101100001010000111001000101010000001111001011000011010; end
            14'd2250 : begin out <= 64'b0010011111011111001010001110011000101001011110011010101000101101; end
            14'd2251 : begin out <= 64'b0010101110110111101001100011010100101010100000110010101010000011; end
            14'd2252 : begin out <= 64'b0010100111100100101001100010011100101011001000100010011010110001; end
            14'd2253 : begin out <= 64'b1010000011000101101010100011010000101000100010111010100010110110; end
            14'd2254 : begin out <= 64'b1001111001110101101010100001110110101000111011010010000000111111; end
            14'd2255 : begin out <= 64'b0001101000101111001010100011000010101001110111111010100110101100; end
            14'd2256 : begin out <= 64'b1010000101010111100111011110101110101000100101110010101101101101; end
            14'd2257 : begin out <= 64'b0010101101110101100100100110010110101011011110010010101110111110; end
            14'd2258 : begin out <= 64'b0010011000111000001000111101110010100100000110100010101101110011; end
            14'd2259 : begin out <= 64'b1010011110100001001010001110110110010110000110110010100011111101; end
            14'd2260 : begin out <= 64'b0010101011111100001000001010001100100100001010111010100000100000; end
            14'd2261 : begin out <= 64'b1001110110010010101010110000011110100110100010101010011101110111; end
            14'd2262 : begin out <= 64'b1010101010111100001001100101000110101011011100010010011001110110; end
            14'd2263 : begin out <= 64'b1010010100011011101010011100100110100111111110000010010011101010; end
            14'd2264 : begin out <= 64'b1010010011101101101010110000101010100001101011110010101001100101; end
            14'd2265 : begin out <= 64'b0010101110110111101010001000101000010011110011101010101100001010; end
            14'd2266 : begin out <= 64'b1010101110010011101010011011001110100110100100111001010011100111; end
            14'd2267 : begin out <= 64'b0010101100111011100100011011000100100111011111110010100111010111; end
            14'd2268 : begin out <= 64'b0001101011101100101010101010011000101011010110101010101000101011; end
            14'd2269 : begin out <= 64'b1010100101100011001010000000000110101000011111101010100001000010; end
            14'd2270 : begin out <= 64'b1010100100010111001010110111110110100101101110010010101101001001; end
            14'd2271 : begin out <= 64'b1000001010101100001000001110111010100100011001101001111110110001; end
            14'd2272 : begin out <= 64'b1010100111010000101010000011101010101011011111100010000110001100; end
            14'd2273 : begin out <= 64'b0001101110000001001000111110100110101011101110100010010011101100; end
            14'd2274 : begin out <= 64'b1010100111000000101010100101010100100100010100110010100110100011; end
            14'd2275 : begin out <= 64'b0010101111110010001010011010101000100111011011110010011000011110; end
            14'd2276 : begin out <= 64'b1010101100111111001010101111110100101011010000100010011101100111; end
            14'd2277 : begin out <= 64'b1010101101010110001001111110100100101011010111001000110010111101; end
            14'd2278 : begin out <= 64'b1010100011011101101001010001011110100100000110101010100011100101; end
            14'd2279 : begin out <= 64'b0001100001010000101010010100000100100111101111101010101101000001; end
            14'd2280 : begin out <= 64'b1010101000100101101010011001011100101001010101011010010001110010; end
            14'd2281 : begin out <= 64'b1010101010101101001001111110100010101011001110101001110010101001; end
            14'd2282 : begin out <= 64'b0010101111111111001001101100011110011110110110100010100011101101; end
            14'd2283 : begin out <= 64'b0010011011010110001001110010111100100011000100001010010101110001; end
            14'd2284 : begin out <= 64'b1010101010100011101010011001111100101010100011000010011101000101; end
            14'd2285 : begin out <= 64'b0010101101101110100100010100111010101011010010111010100111101011; end
            14'd2286 : begin out <= 64'b0010100010101111001001110100100000011110010111001010100001010011; end
            14'd2287 : begin out <= 64'b1010011111111101001001100001100100100101100000010010100100011111; end
            14'd2288 : begin out <= 64'b0010010001001001101010110010101110101010000111010010100000110101; end
            14'd2289 : begin out <= 64'b1010101000111001000111011101011100101001001101101010100011011111; end
            14'd2290 : begin out <= 64'b0000100111100011101010101010101110100010111011101010010101000011; end
            14'd2291 : begin out <= 64'b1010011111001100101010100101101110101010001101011010100111001010; end
            14'd2292 : begin out <= 64'b1010100111000111001010101100111100100110000100011010101001111010; end
            14'd2293 : begin out <= 64'b1010101100101111000111011001100110100100000001010010011011110001; end
            14'd2294 : begin out <= 64'b0010001000000000001010100010010100101011011011101010101100001000; end
            14'd2295 : begin out <= 64'b1010000110001010101000010001101010100011011010101010101111000101; end
            14'd2296 : begin out <= 64'b1010000101101100101001011100011100101011101000000010100110110100; end
            14'd2297 : begin out <= 64'b1010010111111001001010111011101110101010000001100010011110100010; end
            14'd2298 : begin out <= 64'b1010100000001010001010101101001110100101100101001010101001100111; end
            14'd2299 : begin out <= 64'b0001100101110110101010000100000110011001000001001010001011100100; end
            14'd2300 : begin out <= 64'b1010000001000011001010100110011110100100110011110010100101011110; end
            14'd2301 : begin out <= 64'b0010000110000110101010010011110110100111010000100010101010000010; end
            14'd2302 : begin out <= 64'b0010100111110011001000001110010100100110001001110010100100001001; end
            14'd2303 : begin out <= 64'b1001100101111000001010111000011000010111011011101010100010001001; end
            14'd2304 : begin out <= 64'b1010010101010101100100011110101000011111110101010010100011110111; end
            14'd2305 : begin out <= 64'b1010101100000111101001001110011100100101101001100010010001010001; end
            14'd2306 : begin out <= 64'b1010010111110111001010110111101100100101111001000010101000101000; end
            14'd2307 : begin out <= 64'b0010101001100000101010010001101000101001001011110010011001110001; end
            14'd2308 : begin out <= 64'b1010010101010000101010101101100100101000001101000010001111101001; end
            14'd2309 : begin out <= 64'b1010100011100100001001110111100110101011001100100001110010000100; end
            14'd2310 : begin out <= 64'b0010101111010001001010001001010000101001100011001010101000111000; end
            14'd2311 : begin out <= 64'b1010100000011111101010000101111100101010101100111001111110000111; end
            14'd2312 : begin out <= 64'b0001111101011000101000011010000100100101111111110010010011100111; end
            14'd2313 : begin out <= 64'b1010100111111000101010101111111110101010100011100010011111010000; end
            14'd2314 : begin out <= 64'b1010010101101001001010110110001110100110110100101010101110001101; end
            14'd2315 : begin out <= 64'b0010100000011000001010100100000100101010100111111010100101111100; end
            14'd2316 : begin out <= 64'b1010110000000001000111110010010100011110000011111010100011001001; end
            14'd2317 : begin out <= 64'b1010100111100101001010010011101010100110111101000010011000110101; end
            14'd2318 : begin out <= 64'b1010001001101110001010001110010000101010110101101010010011100111; end
            14'd2319 : begin out <= 64'b0010100111001011101001101111001000100110111011001010010001110110; end
            14'd2320 : begin out <= 64'b0010010001011101101010101110111010101000101000010001110010110110; end
            14'd2321 : begin out <= 64'b0001111000001101101001111000011100010011000110111010101001000101; end
            14'd2322 : begin out <= 64'b1010101010101001001010000011011110101001101011110010100111110111; end
            14'd2323 : begin out <= 64'b1010011110000011000110111011100110101000100101001010100010100000; end
            14'd2324 : begin out <= 64'b0001111011001110101010011111100010101000000100001010101100110110; end
            14'd2325 : begin out <= 64'b1010101001111110001010111010010110101000101001000001001010010000; end
            14'd2326 : begin out <= 64'b1010101000000001001010101011000110100010110101111010100000101000; end
            14'd2327 : begin out <= 64'b0001110000111111001001010011101110101001101111101000010011000111; end
            14'd2328 : begin out <= 64'b0010101110010011101010011101110010101001001111101010100101000000; end
            14'd2329 : begin out <= 64'b0001110010111111001000111000110100100011010111001010001111101000; end
            14'd2330 : begin out <= 64'b1010011000010001001010110001001100101011111101001010101110000001; end
            14'd2331 : begin out <= 64'b0010100001110101001000110111110000101000110001011010011010010011; end
            14'd2332 : begin out <= 64'b0010011101011011101010001010101100100111011111000001111010101011; end
            14'd2333 : begin out <= 64'b0010101111011100100111010000010000100110111101000010011001001011; end
            14'd2334 : begin out <= 64'b0010101100011100101010100000110110100100100101101010101000110110; end
            14'd2335 : begin out <= 64'b0010000111000100001001110001010010100111001111100010100111010110; end
            14'd2336 : begin out <= 64'b0010011110101000001001010100100010101001011100100010100000100001; end
            14'd2337 : begin out <= 64'b1010000110101011001010110111101100101001100000011010100000010010; end
            14'd2338 : begin out <= 64'b1010101000011000001010000010001110100111001110010010011010100110; end
            14'd2339 : begin out <= 64'b1010100111011110101000001000000010101010111011001010001011100001; end
            14'd2340 : begin out <= 64'b1010101000001011001001011101100110100001000011101010101000110100; end
            14'd2341 : begin out <= 64'b0001100110101101001000100011000000100100010000000010100100011110; end
            14'd2342 : begin out <= 64'b0010101111000001001010101101111010101010110000100010100101110011; end
            14'd2343 : begin out <= 64'b0010100111111000001010011101000010101011101101110010100011001111; end
            14'd2344 : begin out <= 64'b1010101001001100001010111100100000101001000000100001110000101101; end
            14'd2345 : begin out <= 64'b0010010110010111001000010110100000010000101011010010001100011110; end
            14'd2346 : begin out <= 64'b1010010111000111001010000010110010011010101100000010011110001001; end
            14'd2347 : begin out <= 64'b0010010010101001001010101110011110101011011100101010011110100100; end
            14'd2348 : begin out <= 64'b1010101011100110101010000110011010100111000010000010110001000110; end
            14'd2349 : begin out <= 64'b1010101000000010101010101011111010100101010011100010011010011010; end
            14'd2350 : begin out <= 64'b1010100101110011001001011000101010100111100110101010001001100111; end
            14'd2351 : begin out <= 64'b1010100100111100001000110110011010101010110101100001101000111111; end
            14'd2352 : begin out <= 64'b1001111101011111101001010101000110100000010001001010101111110101; end
            14'd2353 : begin out <= 64'b0010101110101111001010011010010100011001011011100010000100101101; end
            14'd2354 : begin out <= 64'b1010010000001001101010111100111100101011110110011010101111011111; end
            14'd2355 : begin out <= 64'b0001010111001001001010001111011110100100110111010010101000000101; end
            14'd2356 : begin out <= 64'b1010010000100111001000000000001010100111011001111001100010110011; end
            14'd2357 : begin out <= 64'b0010100001110001101010011010010100100100010001110010010001011001; end
            14'd2358 : begin out <= 64'b1010011011100000001010111100101000100111011001000010101011001111; end
            14'd2359 : begin out <= 64'b1010011010011011101010001111010010101000110110000010100111100110; end
            14'd2360 : begin out <= 64'b0010101000001100001010011100010000011101000001011010101110011000; end
            14'd2361 : begin out <= 64'b0010101000010000001001110111011100101000111000001010100000111000; end
            14'd2362 : begin out <= 64'b0010101101101101101010110001001110011101101000000010011000101101; end
            14'd2363 : begin out <= 64'b0010011010100100000110100010001010100001110100010010100011000100; end
            14'd2364 : begin out <= 64'b0010000100110010101010111111111110101010111011111010110000001100; end
            14'd2365 : begin out <= 64'b1010101110010100001001111100010010100011011111001010100011001100; end
            14'd2366 : begin out <= 64'b0010101010110110101010010101101010100101111000011010010011011100; end
            14'd2367 : begin out <= 64'b1010011000111110001010000000011010101001101010110010100011111010; end
            14'd2368 : begin out <= 64'b1001110111010111101001010111111010011110101010101010010110110100; end
            14'd2369 : begin out <= 64'b1001111111001110101001001101011000100111010111000010011000010001; end
            14'd2370 : begin out <= 64'b0010101001001110101010001001101010101001000100111010011101010000; end
            14'd2371 : begin out <= 64'b0010010000010111101010010010000000101011110101001001011000010010; end
            14'd2372 : begin out <= 64'b1010100110000111001010101000110110101011110100001010000100010001; end
            14'd2373 : begin out <= 64'b0010101011111110001001101011000100101001110111011001000110101001; end
            14'd2374 : begin out <= 64'b0010011110110110001010100010111100101011010000111010000110001001; end
            14'd2375 : begin out <= 64'b0001101011100111101001001100001000100000101111111010011100101101; end
            14'd2376 : begin out <= 64'b0010010111100000101001101010101110101010010001110010101000110000; end
            14'd2377 : begin out <= 64'b0010010101110000101001001110011000100111110101001010100110011010; end
            14'd2378 : begin out <= 64'b0010011100010011001001010010101010101001110100111010010010010010; end
            14'd2379 : begin out <= 64'b0010100001001111001001001100000010101011010101101010100100110011; end
            14'd2380 : begin out <= 64'b0010001010110110000101100001000010101011110000010010101001110011; end
            14'd2381 : begin out <= 64'b0010011010001001001000101001101000101001001111011010100000101001; end
            14'd2382 : begin out <= 64'b0010000110010010001010111100010000100001010100111010100010001110; end
            14'd2383 : begin out <= 64'b0010100011100111101000010100100110101000100111001010100110100101; end
            14'd2384 : begin out <= 64'b1010100110101101101010110110100010101010000011010010000100010111; end
            14'd2385 : begin out <= 64'b1010000101100101101010101011011110100110001010000010011111111101; end
            14'd2386 : begin out <= 64'b0001111101111100101001111101010110100011111010100001100110101001; end
            14'd2387 : begin out <= 64'b1010100000011110100110111110101000101000110101011001110111100010; end
            14'd2388 : begin out <= 64'b0010011011000100101010001101101100100000001000110010100111111111; end
            14'd2389 : begin out <= 64'b1010010110101011001010111001000010100011011111101010010011001010; end
            14'd2390 : begin out <= 64'b0010101011100111101000000010100010100100100100110010001100001000; end
            14'd2391 : begin out <= 64'b1010010110010000000111010010010110010101101011010010011010000011; end
            14'd2392 : begin out <= 64'b0010100001101001001001010001100110100010011100010010101100000100; end
            14'd2393 : begin out <= 64'b1001110110001101101010010000010100101001000100111010101110001010; end
            14'd2394 : begin out <= 64'b1001111111001010001001011101111110011100001100110010011000110010; end
            14'd2395 : begin out <= 64'b0010100110011111001010110101111000101000100111111010010010011000; end
            14'd2396 : begin out <= 64'b1010000101110110000110001101010100011110010101101001111111111010; end
            14'd2397 : begin out <= 64'b0010101110010111001010011001101100100011000000010010100000101011; end
            14'd2398 : begin out <= 64'b0010011111011001101010001100100100100101010110100010001011001101; end
            14'd2399 : begin out <= 64'b1010100001100000001010110100010010100100110100101010101011111110; end
            14'd2400 : begin out <= 64'b1001101101100100001010011110100000101000111110001010011111111000; end
            14'd2401 : begin out <= 64'b1001111010011001101001100101001100101000110110111010101101001111; end
            14'd2402 : begin out <= 64'b0001010000011101101001001101110000011111111010110010101000000000; end
            14'd2403 : begin out <= 64'b0001110011010010101000101010010110100011011101100010011101001010; end
            14'd2404 : begin out <= 64'b1010101111101111001001100100000100101000001010011010000101100111; end
            14'd2405 : begin out <= 64'b0010100100000111001010110010110000101010110101110010011011111001; end
            14'd2406 : begin out <= 64'b0010000100100000101001101101000010101000101101000010101001111011; end
            14'd2407 : begin out <= 64'b1010100111101101001010110111001010100111101110111010010010001010; end
            14'd2408 : begin out <= 64'b0010011101000000001010111001101010011101111011001010011001110100; end
            14'd2409 : begin out <= 64'b1010101110110001001010111100011000101010111111000010010111010010; end
            14'd2410 : begin out <= 64'b1010100010100110100011100010110110100101111110000010100000001011; end
            14'd2411 : begin out <= 64'b1010011001101111001010101101101000100100001100000010010101011011; end
            14'd2412 : begin out <= 64'b0010011010011111101001111111011100100100001101111010101001101110; end
            14'd2413 : begin out <= 64'b1010011101100101001010011001010100101011011010101001100100111000; end
            14'd2414 : begin out <= 64'b0010100100110000101010011001010110100001110100011010011001111001; end
            14'd2415 : begin out <= 64'b1010100010111001001010000100100000101000111000000010100011100111; end
            14'd2416 : begin out <= 64'b0010100010011001001001111000001100101010110000100010100010010010; end
            14'd2417 : begin out <= 64'b0010000011101101001001100110101010100111000101011010011010101110; end
            14'd2418 : begin out <= 64'b1010101011101011001010010001011100100011110011101010100101110110; end
            14'd2419 : begin out <= 64'b0010010111010001100000011111111100011100110111110010100110001010; end
            14'd2420 : begin out <= 64'b0010100001110101100100010101010110100000111101101010100110110010; end
            14'd2421 : begin out <= 64'b0010010010001000001001101101010110100011111010010010100011110001; end
            14'd2422 : begin out <= 64'b1010100001100110001010010110011000100101111111110010010101001010; end
            14'd2423 : begin out <= 64'b0001000111000000001010100101111000101000111101000010100110111001; end
            14'd2424 : begin out <= 64'b0010100011001111101010000100100010101000010010101001110010001111; end
            14'd2425 : begin out <= 64'b0010101000100101101010000010111000101011010000100010011001001101; end
            14'd2426 : begin out <= 64'b0010101000111100001001010000100100101100000000101010100101011101; end
            14'd2427 : begin out <= 64'b1010010100111111001010011000001000101010101000100001000100100100; end
            14'd2428 : begin out <= 64'b1010101101111000001001100111000000010111110010101010010100010000; end
            14'd2429 : begin out <= 64'b0010011001011001101010000011111100100111110100001010100011000010; end
            14'd2430 : begin out <= 64'b0010100110010100001001101010100000101001101100110010101000000100; end
            14'd2431 : begin out <= 64'b0010100011101011001010011111101100101001110011000001110111111001; end
            14'd2432 : begin out <= 64'b1010101000111101000111100010000110101010100100101010101001110101; end
            14'd2433 : begin out <= 64'b0010100100100001001010001110001110100100110101100010001000011000; end
            14'd2434 : begin out <= 64'b1010101000100110101000101010101000101011110011011010101101010001; end
            14'd2435 : begin out <= 64'b1001001010100000001010011100000100101010010111110010010000010010; end
            14'd2436 : begin out <= 64'b1001111001000101001010000101000010100110101100001001110010111111; end
            14'd2437 : begin out <= 64'b0010001101001000001010001010000100100011000011111010100100000101; end
            14'd2438 : begin out <= 64'b0010101101001100001010110101111000101010000111001010010010011101; end
            14'd2439 : begin out <= 64'b0010101001111110101010000000111100100100110100011010011111000000; end
            14'd2440 : begin out <= 64'b1010100001000110100101110000111100100001010101100010000110100110; end
            14'd2441 : begin out <= 64'b0010010001011010101000000110110110100001100001011010100110100001; end
            14'd2442 : begin out <= 64'b1001111001011110001010000001110010100011011111110010001110110110; end
            14'd2443 : begin out <= 64'b0010100110001001001001101001100100010000110010110010101100100101; end
            14'd2444 : begin out <= 64'b0010100111101111101010101000000110101000100101111010100101011101; end
            14'd2445 : begin out <= 64'b0010010110011010100110000101010100100111111001111010100011101011; end
            14'd2446 : begin out <= 64'b1010100010111110101011000001101110100100011001111010010100110110; end
            14'd2447 : begin out <= 64'b1010101011110001101000111001000000101001111110111010011011101010; end
            14'd2448 : begin out <= 64'b1010010100101100001000000001001000101001001000100010101101111001; end
            14'd2449 : begin out <= 64'b0010011010100111101011000000100100101000010010000010101101101011; end
            14'd2450 : begin out <= 64'b1010010101001010101010011001011100011101101111011010000001100010; end
            14'd2451 : begin out <= 64'b0010100010101101001000010001101100011001110100101001110110010100; end
            14'd2452 : begin out <= 64'b1010101010111011001010001001101000101000111101011010010100111011; end
            14'd2453 : begin out <= 64'b0010011101001010001010110010101000011100111111101010100111001110; end
            14'd2454 : begin out <= 64'b0001010011111010001001011011000100101011110001000010011111110001; end
            14'd2455 : begin out <= 64'b1010100011111111100111000001101000101001000110101010000110101001; end
            14'd2456 : begin out <= 64'b1010101111001000101010011111101110100100111110000010101010000010; end
            14'd2457 : begin out <= 64'b1010100100101000101010001001000100101011010101011001100001010011; end
            14'd2458 : begin out <= 64'b0010100001000101001010110000000110100001011011001010011011100110; end
            14'd2459 : begin out <= 64'b1010000011000001101001110000001110100110111011101010101001110111; end
            14'd2460 : begin out <= 64'b1010101101001010100100100011101000101011000101000010010001010000; end
            14'd2461 : begin out <= 64'b1010100111101001001010100011110000100000001001100010010101110110; end
            14'd2462 : begin out <= 64'b1010010001111111101010100000101010100011100101101010100111010101; end
            14'd2463 : begin out <= 64'b0010101110100000001001101101110100100111110111001010101110011111; end
            14'd2464 : begin out <= 64'b0001100011110111001001110001111110100101010101111010001000110000; end
            14'd2465 : begin out <= 64'b0001111010000101001010110011000100101001010111001010100110001110; end
            14'd2466 : begin out <= 64'b0010101100100100001001111010001100101011011111000001101001110111; end
            14'd2467 : begin out <= 64'b1010010010011001001010001100001010100011011101001010001001001001; end
            14'd2468 : begin out <= 64'b1010100001111111000000011110100000101001001100001001001001111011; end
            14'd2469 : begin out <= 64'b1010101100110001101010100001001010010110110110100010000100100110; end
            14'd2470 : begin out <= 64'b1001101000101001101010101010101100011101101000110010100000011100; end
            14'd2471 : begin out <= 64'b0010101010010011101010101110011010101001010010110010100100000111; end
            14'd2472 : begin out <= 64'b1010010101001100101000111010111100101010000111111010011100000111; end
            14'd2473 : begin out <= 64'b0010101100000011101010001110010100101010110111111001111000001000; end
            14'd2474 : begin out <= 64'b1010010111010000001010001001000010100101100101010010100100000001; end
            14'd2475 : begin out <= 64'b0010101010000111001010111101101110011111010110001010001011111110; end
            14'd2476 : begin out <= 64'b1001101100110001001010100110010100101000100100000010011100100111; end
            14'd2477 : begin out <= 64'b0010100001110100001000000010001110101011011001001010101111100110; end
            14'd2478 : begin out <= 64'b0010100101101010101010110001001100100110001001011010011000010111; end
            14'd2479 : begin out <= 64'b1010010001011010000111111000001110101011000100000001110001001010; end
            14'd2480 : begin out <= 64'b1001111111111101001000010101011110100101111110000010011111001101; end
            14'd2481 : begin out <= 64'b1010100001100101101010000001101100101001000011111010100000110101; end
            14'd2482 : begin out <= 64'b0010011011000100000110100011001110101001111111000010101010010000; end
            14'd2483 : begin out <= 64'b1010101101110000000111001000110010100111100110001010011010100010; end
            14'd2484 : begin out <= 64'b1010100101100101101010001001100110100010001110101010100011110101; end
            14'd2485 : begin out <= 64'b0010100111101110001010100111100000101000000100000010101101011011; end
            14'd2486 : begin out <= 64'b0010101101111001100101010111101100100100001100001010100111001011; end
            14'd2487 : begin out <= 64'b1010100011001111001010011000101010011101000010101010101111001011; end
            14'd2488 : begin out <= 64'b1010011010011011001001100001000110101001010110000001100110001111; end
            14'd2489 : begin out <= 64'b1010101100000001001001010001001100101000000010100010101001001001; end
            14'd2490 : begin out <= 64'b1010010110100101101010001001110110101011010000010010101001110001; end
            14'd2491 : begin out <= 64'b0010011101110110001010100010101000011010100011111010010001011011; end
            14'd2492 : begin out <= 64'b1001000110000011101010001011000000101000010101000010001111011110; end
            14'd2493 : begin out <= 64'b0010010111100010101001101011101000101000100101110010100111110100; end
            14'd2494 : begin out <= 64'b1001100111011101101010101111010010100111010110101010101001110100; end
            14'd2495 : begin out <= 64'b0010101011010110101010101001000010100100001010110010100100011011; end
            14'd2496 : begin out <= 64'b1010011010110111001011000000000110101010001111010010100101010110; end
            14'd2497 : begin out <= 64'b0010100101101000101010110111101000101010000001010010100001101111; end
            14'd2498 : begin out <= 64'b0010101101001001101000000101010100100101111100000010001110000111; end
            14'd2499 : begin out <= 64'b0010000010000110001010100100110100101001110010110010100011010001; end
            14'd2500 : begin out <= 64'b1010010110011000001001010100000100011110110011111001100110110001; end
            14'd2501 : begin out <= 64'b0010011110110011001001000101110100101000111000011010001000010100; end
            14'd2502 : begin out <= 64'b1010001110001011101000000110000100101011000110011010101110101110; end
            14'd2503 : begin out <= 64'b0010100011110011001001001011001000100111010001100010100111100001; end
            14'd2504 : begin out <= 64'b1010100111010000101010101000000010101001010000001010100100111001; end
            14'd2505 : begin out <= 64'b1010100100010101000110111110101100100111010011001010011001100100; end
            14'd2506 : begin out <= 64'b0010101011111111101010001101101000100101000111111010101011101111; end
            14'd2507 : begin out <= 64'b1010101100000100101000100101010100101000101110111010010001011000; end
            14'd2508 : begin out <= 64'b1010101110100111101010100101111010100101101111000010101101010000; end
            14'd2509 : begin out <= 64'b1010001011000011001001100010100010100110100001111010010011100100; end
            14'd2510 : begin out <= 64'b1010101010111011001010101110011110100111010001001010010110110111; end
            14'd2511 : begin out <= 64'b1010101101010011001010011110011110101001001000110010101010000101; end
            14'd2512 : begin out <= 64'b1001110011000000101010011101100100101000000110111010011100101010; end
            14'd2513 : begin out <= 64'b1010100001110011100110010111101010101000000101110010101000100110; end
            14'd2514 : begin out <= 64'b0010101111011111001010001010001110100100110000111010100110000100; end
            14'd2515 : begin out <= 64'b1010101000001101101001010001101100011001001110110010011111011111; end
            14'd2516 : begin out <= 64'b0010101100101011001001010111101010100000100111100010101011100010; end
            14'd2517 : begin out <= 64'b1010100010101110101001000100010110011010101110000010100101011001; end
            14'd2518 : begin out <= 64'b0010100111010101001010011111011010011111000001100010101001001110; end
            14'd2519 : begin out <= 64'b0010001111100010101010001010100100100010000001100010101011000110; end
            14'd2520 : begin out <= 64'b0010101011100100100111100001110110101001100110110010000001001010; end
            14'd2521 : begin out <= 64'b0010101100111110001010110000011100100101011001110010100101001001; end
            14'd2522 : begin out <= 64'b1010011111000001100110001111000110001001010101010010101011110111; end
            14'd2523 : begin out <= 64'b1010000111010011000111000001001010101000111000100010000000100101; end
            14'd2524 : begin out <= 64'b0010001000000000101010000101010010011110101001010010101110100100; end
            14'd2525 : begin out <= 64'b0010001011101000101010100001110110100100111100110010000001101110; end
            14'd2526 : begin out <= 64'b1010101010010101101010001011101110011011101001011010101111101110; end
            14'd2527 : begin out <= 64'b1001111110110100100110111000100010100101000000011001111000001001; end
            14'd2528 : begin out <= 64'b0010010000010110001010000111100000100100110001001010000100110110; end
            14'd2529 : begin out <= 64'b1010010011110110001010101110011110100110110100010010010110110111; end
            14'd2530 : begin out <= 64'b0010100000100010100111110000111110101000010010100010101111000011; end
            14'd2531 : begin out <= 64'b0010100111101011101001011101100100101000011111010001010100100001; end
            14'd2532 : begin out <= 64'b0010101100110001101001001110100110010101110101111010010110101110; end
            14'd2533 : begin out <= 64'b0010000111010100001001000000100110100110101000111010101101101010; end
            14'd2534 : begin out <= 64'b1001011010010010101000010111100000101001101001001010100110000101; end
            14'd2535 : begin out <= 64'b1001100011011100001010110110010100101010110111010010100111110000; end
            14'd2536 : begin out <= 64'b0010010111111101001000111110101110101011111110100010101010110010; end
            14'd2537 : begin out <= 64'b0010100010100101101010111110010010101010111110001001110111001111; end
            14'd2538 : begin out <= 64'b1010101100011111000110101111011010101000110010100010100100111000; end
            14'd2539 : begin out <= 64'b0010010010001101100111100100010010100001111010001001100010000111; end
            14'd2540 : begin out <= 64'b0010001111100001001010111011010100100000100011010010011001000001; end
            14'd2541 : begin out <= 64'b0010010001001001101010001101010010100000010010110010101100111000; end
            14'd2542 : begin out <= 64'b1000110100000011101010110011100000100100001111011010100001011111; end
            14'd2543 : begin out <= 64'b0010011010100110001010110011111000101000110101101010101100101010; end
            14'd2544 : begin out <= 64'b0010001001111010101010110100100110100101100110100010101011000100; end
            14'd2545 : begin out <= 64'b0010101100010000101010110101111100100111101001110010000101011011; end
            14'd2546 : begin out <= 64'b0010100000111001001010101011001110100111111010011010100110001011; end
            14'd2547 : begin out <= 64'b1010101001000110101001001110101010100000010101001010011001111001; end
            14'd2548 : begin out <= 64'b1001110111111010001010010011010000101011100010000001011001001011; end
            14'd2549 : begin out <= 64'b1001110101100110001001000000100100101010100111001010100100000101; end
            14'd2550 : begin out <= 64'b1010010010001101101010111000101100101000000000001010101000011110; end
            14'd2551 : begin out <= 64'b1010101101010011100111011010111010101010010110100010000001111101; end
            14'd2552 : begin out <= 64'b0010100111001001001001110010011000101011100101111010010011111111; end
            14'd2553 : begin out <= 64'b1010101010111011101010001111001100100001001111010010101011000110; end
            14'd2554 : begin out <= 64'b1010001010110101101000101010011100100111100101010010101111100100; end
            14'd2555 : begin out <= 64'b1001011010001010101001111000001100101001110000000010101111010011; end
            14'd2556 : begin out <= 64'b0010100011100001101000101000101010101000011111111010010000100100; end
            14'd2557 : begin out <= 64'b1010100110101000101001100101010000101001101110101001110111110111; end
            14'd2558 : begin out <= 64'b0010100000000110101001011010101000100001101100111010011001010110; end
            14'd2559 : begin out <= 64'b0010011001101001001000111101101110101000011101101010100000011011; end
            14'd2560 : begin out <= 64'b1010101011110111000111111110101000101001111101001010100001101101; end
            14'd2561 : begin out <= 64'b0010100101011000001010100001111010001001011111111010010001111010; end
            14'd2562 : begin out <= 64'b1010100010011101000110110100001000101011000101010010100000010011; end
            14'd2563 : begin out <= 64'b1010000011001001101000110100011100101010001100011010010100101011; end
            14'd2564 : begin out <= 64'b1010010110100010001000000110100010100111101011011010101000100011; end
            14'd2565 : begin out <= 64'b0010101011010110001001101000011110100111110100111010101001000101; end
            14'd2566 : begin out <= 64'b1010101010100011100100001000101110100011111100110010000001000001; end
            14'd2567 : begin out <= 64'b0010100111000111101010100110001010100101010000010010011110010110; end
            14'd2568 : begin out <= 64'b1010101010110000001010010010110010100111010011101010000110111001; end
            14'd2569 : begin out <= 64'b0010100010100101001010010111100110100100001101000010101001100000; end
            14'd2570 : begin out <= 64'b0010101101101100001011000001100000100011111100111010011101111010; end
            14'd2571 : begin out <= 64'b0001001001010100001010100011010100100000110010011010100111010110; end
            14'd2572 : begin out <= 64'b1010100000111000101010011011111000011111100100011010010011001101; end
            14'd2573 : begin out <= 64'b0010011100111001100111000101101000101000010010011010000011111110; end
            14'd2574 : begin out <= 64'b0010101000000010000110100010111000101010111000001010011110101100; end
            14'd2575 : begin out <= 64'b1010011100101111101000101001111110100010111110000010011000000110; end
            14'd2576 : begin out <= 64'b1010010000100101001010101111001000100110001101001010100111110111; end
            14'd2577 : begin out <= 64'b0010000100101000101010000001000010011001001111001010100000011110; end
            14'd2578 : begin out <= 64'b0010100100100010101010010111010110101001000111100001110100001000; end
            14'd2579 : begin out <= 64'b1010101011100001101000000111001100010011100110100010101001110000; end
            14'd2580 : begin out <= 64'b0010101011100110101010010110000010011100001111001010011100101101; end
            14'd2581 : begin out <= 64'b1010001010010110001001010111101100101010101110010001110001100111; end
            14'd2582 : begin out <= 64'b1001111101000001101010100111011010100001001000101010010101110011; end
            14'd2583 : begin out <= 64'b0010100001011000101000010010010100101011100100001010101010010000; end
            14'd2584 : begin out <= 64'b0010100010111010001010001001000100011110011101110010100110001000; end
            14'd2585 : begin out <= 64'b1010101101100101101010110001111010100011100110111010011010010101; end
            14'd2586 : begin out <= 64'b1010100001111100001010011100100100100110011000100010101100110010; end
            14'd2587 : begin out <= 64'b1010101011000000100111011000111100101001010101101010000000100001; end
            14'd2588 : begin out <= 64'b1001100011000100101000111011001000101010100110111010101110001000; end
            14'd2589 : begin out <= 64'b0010100100010011101010000000000110011101101110000010100101010100; end
            14'd2590 : begin out <= 64'b1010010010111100001011000000110010011111110010001010100001100010; end
            14'd2591 : begin out <= 64'b1001111010100110101000010010010000101001010100100010101011011100; end
            14'd2592 : begin out <= 64'b0010000010111011101010101001010100011110001000111010010100111101; end
            14'd2593 : begin out <= 64'b1010000110000110101000001100111100101010010001100010000011111010; end
            14'd2594 : begin out <= 64'b0010100111111101001010001010100100101001011111100010100101010011; end
            14'd2595 : begin out <= 64'b1010100100011111000111011100110000100001100000011001110100000011; end
            14'd2596 : begin out <= 64'b0010001001011001100101100011001000101011001101001010100100111000; end
            14'd2597 : begin out <= 64'b1010010111100001001010110010100100101001101000100010011101010101; end
            14'd2598 : begin out <= 64'b0001101110001001101010001111000100101000101001001010100010001101; end
            14'd2599 : begin out <= 64'b1010000010000111001000010110000000101011010011011010101000110101; end
            14'd2600 : begin out <= 64'b1001011010111110001001111011000100001110100110011010101000110001; end
            14'd2601 : begin out <= 64'b0010101011100101101001111010001000101001001101101010101011101010; end
            14'd2602 : begin out <= 64'b1010011101101100101010111010010010100100001111010010101011111100; end
            14'd2603 : begin out <= 64'b0010001111110110101000111001100010100100100110011010100101111101; end
            14'd2604 : begin out <= 64'b0010100001110100101010101011010110101001101111010010000101010100; end
            14'd2605 : begin out <= 64'b0010010011011010001001110101101000100100010011100010100010000001; end
            14'd2606 : begin out <= 64'b1010100111111110101010101110100110011011100010101010010110110111; end
            14'd2607 : begin out <= 64'b1010000110100110101010110000110000100100001000010001101110001100; end
            14'd2608 : begin out <= 64'b0001100000101000101010001011100110101011000111011010101111110111; end
            14'd2609 : begin out <= 64'b0010100101001000001010101110000000101010000100000010101011101000; end
            14'd2610 : begin out <= 64'b1001110111101100001001000001101000101000111101110010100101010111; end
            14'd2611 : begin out <= 64'b0010100010110110101001010100011010100011101000110010100001011111; end
            14'd2612 : begin out <= 64'b0010101101001110001000010011011100010011100010111010100100010000; end
            14'd2613 : begin out <= 64'b1010101110000000101010100100011100101010110100110010100100100000; end
            14'd2614 : begin out <= 64'b1010100111000001101000100110011110100101111001101010101110110010; end
            14'd2615 : begin out <= 64'b0010100110001001001011000000101010100101100011110010010111011101; end
            14'd2616 : begin out <= 64'b1010101001011000001010011101011000101001001100000010100011010111; end
            14'd2617 : begin out <= 64'b0010100011100010001010111110110100101010110101100010100111011001; end
            14'd2618 : begin out <= 64'b1001100101101110001001001000111000100111101001000010100000011000; end
            14'd2619 : begin out <= 64'b1010101110001101001010010011101000101011000101111001111111111011; end
            14'd2620 : begin out <= 64'b1010001101110100000111011001101010101000001010111010101000000000; end
            14'd2621 : begin out <= 64'b0010101000110110001001001001101100101010011001001010100011011010; end
            14'd2622 : begin out <= 64'b1010100111100001001010010000111000101010011010110010011010100101; end
            14'd2623 : begin out <= 64'b0010100010101000001001001111011110100001101101000010000010111100; end
            14'd2624 : begin out <= 64'b0010100110001110101000100100001000100000011110111001010111100011; end
            14'd2625 : begin out <= 64'b1010100101111110001011000011000000100111010100011010000001011010; end
            14'd2626 : begin out <= 64'b0010001001111001001001110101010000100100000011101010100010101011; end
            14'd2627 : begin out <= 64'b1010011010011100001010010110100110100100010011000010010001011101; end
            14'd2628 : begin out <= 64'b0010100100011100101001111001000110100000110010111010010110100101; end
            14'd2629 : begin out <= 64'b0010010110101101001001011111100000100011100011110010000101011010; end
            14'd2630 : begin out <= 64'b0010100101111110101010011110111110010110101011001010101100111001; end
            14'd2631 : begin out <= 64'b1010100110101010101010110111101100100011000011001001101110110000; end
            14'd2632 : begin out <= 64'b1010100100111100101010011110011100011101001010101010010111101101; end
            14'd2633 : begin out <= 64'b0010010110101010001010110100010100101001001110101010101010010110; end
            14'd2634 : begin out <= 64'b1010001010000001101010111011001000100010111001111010100011000001; end
            14'd2635 : begin out <= 64'b0010101110010000001010000011010010101010100010110010010000100101; end
            14'd2636 : begin out <= 64'b1010011100101010101010110010001110101011110111000010101001100100; end
            14'd2637 : begin out <= 64'b0001011101101000100110001000110010101011100100110010101011110001; end
            14'd2638 : begin out <= 64'b1010001000110000100101100100100010100110111000110010011110110011; end
            14'd2639 : begin out <= 64'b1010010100001110001010101001010000100111100110110010110000000101; end
            14'd2640 : begin out <= 64'b0010011001010011000011101011110110100011110011001010010010101110; end
            14'd2641 : begin out <= 64'b1010101011011110101001010010101000100101100011000010010001000100; end
            14'd2642 : begin out <= 64'b1010100101001101100101011010111000101011110110100010011011101111; end
            14'd2643 : begin out <= 64'b1010101010110010101010000000011100101010110101010010010101000011; end
            14'd2644 : begin out <= 64'b0010010000111011101010110100100110011110111101110010101000000001; end
            14'd2645 : begin out <= 64'b1010100111110100100110001001001000101010111110100010101011011010; end
            14'd2646 : begin out <= 64'b1010101111001101000111111101001000101001001000101001110000101110; end
            14'd2647 : begin out <= 64'b0001011000000000101010110011110000011010100010101010100010111110; end
            14'd2648 : begin out <= 64'b0010011001101111001010110011010010101000111111011010101001111011; end
            14'd2649 : begin out <= 64'b0010011110111110001010001010110110011100011011011010001110001111; end
            14'd2650 : begin out <= 64'b0010010011110111001000011010010100101001001110011010011100101101; end
            14'd2651 : begin out <= 64'b1010011100101111101001000111011010011110011000000010011101011000; end
            14'd2652 : begin out <= 64'b1010101011111110100110011111011110101010001100001001110101010010; end
            14'd2653 : begin out <= 64'b0010101001000010001010110101001000101010000111101010100011110101; end
            14'd2654 : begin out <= 64'b1010011001110001000111001101000010100010001001001010101100011000; end
            14'd2655 : begin out <= 64'b0010011001110100101010101011000000100100001110110010101100101010; end
            14'd2656 : begin out <= 64'b0010001011011100000110100011100010101010011011011001111001101001; end
            14'd2657 : begin out <= 64'b1001110001110110101010110101110110100001000011010010101000110110; end
            14'd2658 : begin out <= 64'b1010100110111100001010111000111000101011110000001010000000010111; end
            14'd2659 : begin out <= 64'b0010100111010100101010011001101100101001000100110010100101101000; end
            14'd2660 : begin out <= 64'b0010101110111111001001010010111000100011010110001010101011011000; end
            14'd2661 : begin out <= 64'b1010101101110110100110011001011110011010010000001010100001001101; end
            14'd2662 : begin out <= 64'b0010001111111011000011001110100010101000010011011010101111001001; end
            14'd2663 : begin out <= 64'b0010101100100101101001111111000000101011001011001010101011010011; end
            14'd2664 : begin out <= 64'b1010101001000110001001111000011110100011001101110001110010011001; end
            14'd2665 : begin out <= 64'b0010001100001000001000011011100000101010011111001010101001101000; end
            14'd2666 : begin out <= 64'b0010101101001100101010111010000100100100101110110010000001110011; end
            14'd2667 : begin out <= 64'b1010100100001111001010010010111110101010100101011010101110011001; end
            14'd2668 : begin out <= 64'b0010010111100010001000011111100110100100001010001010101000000000; end
            14'd2669 : begin out <= 64'b1010101111100101101001000010001100100011011110000010101000000111; end
            14'd2670 : begin out <= 64'b0010011100011001001001101010110100101000000011111001101001001001; end
            14'd2671 : begin out <= 64'b0010100101101011001010001111110100100100010010000010110000011000; end
            14'd2672 : begin out <= 64'b1010100111001100001010010111100000100101100101100010100110000011; end
            14'd2673 : begin out <= 64'b1010100111001101101010001000101110100010000000011010010001110010; end
            14'd2674 : begin out <= 64'b1010001001010000001010110010000100011001110000001010010010011101; end
            14'd2675 : begin out <= 64'b1010011101011010001001111010111110101010110101100010011011110100; end
            14'd2676 : begin out <= 64'b0010100110011100001010000011001100100110110100000010100110011011; end
            14'd2677 : begin out <= 64'b0010100101110010000111101111001100101011001110101010100010101111; end
            14'd2678 : begin out <= 64'b0001111100100001101001100100011000100110000101000010011100111001; end
            14'd2679 : begin out <= 64'b0010101100110111001010001101101100100100001011000010011000010110; end
            14'd2680 : begin out <= 64'b0010101111000100101010001110010110100101000110000010001101011100; end
            14'd2681 : begin out <= 64'b1001111101001100001001001111111000100101101010011010010110110101; end
            14'd2682 : begin out <= 64'b0010100000001101001010000010011000100011001001011001110000110010; end
            14'd2683 : begin out <= 64'b0010101101111001101010011001100100100100000111110010100110001011; end
            14'd2684 : begin out <= 64'b0010101100011000100111000110101000011101111001101010100000101011; end
            14'd2685 : begin out <= 64'b1010010010011101101010010000111010101010111110100010101110001001; end
            14'd2686 : begin out <= 64'b1010101010111100001000100010101000011101010011111010011000111111; end
            14'd2687 : begin out <= 64'b0001000000111101001010101101101010100111001111111010010101101011; end
            14'd2688 : begin out <= 64'b1010100111010001101010000000100110101001110100001010011011001111; end
            14'd2689 : begin out <= 64'b1001010111111101001000010101110110100100110101011010100010100110; end
            14'd2690 : begin out <= 64'b0010101001000111001010001101100110101000110000011010100111000110; end
            14'd2691 : begin out <= 64'b1010011101100011101010101011000000100110111110001010101010111001; end
            14'd2692 : begin out <= 64'b0010100010000010000110000100000000101001101011110010011000111100; end
            14'd2693 : begin out <= 64'b0010100110110101001010011010011000100001000100110010011001010100; end
            14'd2694 : begin out <= 64'b0010101000111101001001001000100110101010000111001010011001000101; end
            14'd2695 : begin out <= 64'b0010100111001001101001100110111110100110101001001000000110111010; end
            14'd2696 : begin out <= 64'b1010101100100010001000111101110010101001000011101010100010100011; end
            14'd2697 : begin out <= 64'b1010100000001001101010001000111000101011010110000010011110011110; end
            14'd2698 : begin out <= 64'b1010011111101101001010000010110000100001111000100010010111010111; end
            14'd2699 : begin out <= 64'b0010011001000101101010001011000100101010100000001010010001110100; end
            14'd2700 : begin out <= 64'b1010101100111111000111110111101000100000000011111010100111000101; end
            14'd2701 : begin out <= 64'b1010011100110101101010110001010100100111111110101010010011011000; end
            14'd2702 : begin out <= 64'b0010101111110010101010010101110110100100000101111010100100110000; end
            14'd2703 : begin out <= 64'b0010101010001101001010111010000010101000110110100010101101001011; end
            14'd2704 : begin out <= 64'b1010100001110101001000011110111100101000010001100010100101101011; end
            14'd2705 : begin out <= 64'b1010010011000000001001101111010000011100110001100010010001001110; end
            14'd2706 : begin out <= 64'b1010100101001011101000110010110100101010000110001001111101111001; end
            14'd2707 : begin out <= 64'b0001110001100011001010010100010010100101100010110010101001011101; end
            14'd2708 : begin out <= 64'b1001011100001010101001101011000000101001010011011010101101110101; end
            14'd2709 : begin out <= 64'b0010100101011101101010010001111110101010101110101010010100010110; end
            14'd2710 : begin out <= 64'b1010011011000001101010110101111010101000100000010010100101110000; end
            14'd2711 : begin out <= 64'b1010101101000001001001101101010010101001111001010010100011010101; end
            14'd2712 : begin out <= 64'b0010101101111110101000111100101000101000110010101010101100100001; end
            14'd2713 : begin out <= 64'b1001110100110101001010000011001100100100111000110010101101110000; end
            14'd2714 : begin out <= 64'b0010101001001001101010100011111110100111011011000010010000100001; end
            14'd2715 : begin out <= 64'b0010010111100111001001111100101110100010100000110010010100100111; end
            14'd2716 : begin out <= 64'b1010100110010001001001111010101100101011110100100010101000011001; end
            14'd2717 : begin out <= 64'b0001100100001010001010111000010000101010100011011010101110011110; end
            14'd2718 : begin out <= 64'b0001000010101101101010000000110110101011011100000010101011001000; end
            14'd2719 : begin out <= 64'b0010001000110011001010011011110100100100101111011010101010101011; end
            14'd2720 : begin out <= 64'b0010010100110110101000011011000100101001111100011010100110101110; end
            14'd2721 : begin out <= 64'b0010101000101110101010101111110010100101010101010010101101011111; end
            14'd2722 : begin out <= 64'b0010101010000011101010011110101000101001100110001010011100000011; end
            14'd2723 : begin out <= 64'b1010011111100111101001111010010000100001011010110010100101000000; end
            14'd2724 : begin out <= 64'b0010010110100101001001000101010000100010001001011010011101110010; end
            14'd2725 : begin out <= 64'b1010100110000001101010110000101100101000010111001010100110011101; end
            14'd2726 : begin out <= 64'b1010000100101100101010001001010000101000011001111010101110011101; end
            14'd2727 : begin out <= 64'b0010011000000100001000000000101010101000100001000010000010100110; end
            14'd2728 : begin out <= 64'b1010100000101110001001000001101100011110001111001010100000101100; end
            14'd2729 : begin out <= 64'b0010101100101001001010010011010000100110010000101010000010111000; end
            14'd2730 : begin out <= 64'b1010100101101001001010000000101100101011101010001010101000010000; end
            14'd2731 : begin out <= 64'b0001110001110010001010100010110010101001001000111010011001000100; end
            14'd2732 : begin out <= 64'b1010011001010101101010000100001100011100111001001010101110111011; end
            14'd2733 : begin out <= 64'b1010101011111001001010110010111100101010101101111001110000110010; end
            14'd2734 : begin out <= 64'b0010010001000111100011000000010110010110100011100010011100101101; end
            14'd2735 : begin out <= 64'b1010101110001110101010100010011010010100101110000010011101110000; end
            14'd2736 : begin out <= 64'b1010100001011111100110001110101010100100111010010010010100011011; end
            14'd2737 : begin out <= 64'b1010101000010011101001111100010110100010010100100010011010100110; end
            14'd2738 : begin out <= 64'b0010101100100101001011000000001100100111010000100001111100111100; end
            14'd2739 : begin out <= 64'b0010101101010011001010001101000000101011110101001010010001001000; end
            14'd2740 : begin out <= 64'b0001100001011001100110000010010100101001100110010010101010000110; end
            14'd2741 : begin out <= 64'b0010101010100110001001110111110010101011000110101010011011000110; end
            14'd2742 : begin out <= 64'b0001011000111010101010000100001110101010011110010010101011011101; end
            14'd2743 : begin out <= 64'b0010101010010111001000111000011100101001100010011010101011001110; end
            14'd2744 : begin out <= 64'b0010101010111111001010011101101000100111010000010010011010001001; end
            14'd2745 : begin out <= 64'b0010010011101010001010001100111100100111001100111010011101111100; end
            14'd2746 : begin out <= 64'b1010010110001101100110000011000100101000010101111010010100000110; end
            14'd2747 : begin out <= 64'b1010011110001001101001010011010100100000010010101000100111000011; end
            14'd2748 : begin out <= 64'b1010101011011111001010101101010100100110101011001010100111111101; end
            14'd2749 : begin out <= 64'b1010011001000000001010110000110110011100110000001010101110111111; end
            14'd2750 : begin out <= 64'b1010010101101110001010001001001010101010111101100010100110110100; end
            14'd2751 : begin out <= 64'b0010010011100001101010100001010110011100100000011010100000111000; end
            14'd2752 : begin out <= 64'b0010100010110010101010011110110110101010100100100010100101110011; end
            14'd2753 : begin out <= 64'b1010100010111010001010110110010010011110101001101010101010000000; end
            14'd2754 : begin out <= 64'b0010101111000011001010001100010110100100111111000010100110001000; end
            14'd2755 : begin out <= 64'b0010010111101010101001000111010000101100000011000010100110000101; end
            14'd2756 : begin out <= 64'b0010101101011010101000010001010100100001001101101010100001001111; end
            14'd2757 : begin out <= 64'b0010011111000000101000111001011110011000110111000010100011101101; end
            14'd2758 : begin out <= 64'b1001110100000011001000011010010000101001000000101010101011110110; end
            14'd2759 : begin out <= 64'b0010001100100100101010010111110110101000000000010010101111010110; end
            14'd2760 : begin out <= 64'b1010100010110010101000100010111110100001001100010010000010101001; end
            14'd2761 : begin out <= 64'b0010010111111011101010000000000010101010101101001010011011010100; end
            14'd2762 : begin out <= 64'b0010011100000000001000010101001110101010110010000010011000110001; end
            14'd2763 : begin out <= 64'b0010101111011100101010011010111010101001001011110010100011100011; end
            14'd2764 : begin out <= 64'b0010101000101100001000010101101000011011100100101010100010100100; end
            14'd2765 : begin out <= 64'b0010101111100011001001110100011010100100000101001010000111110001; end
            14'd2766 : begin out <= 64'b0010101100100010001001000011000010101011000100101010100011100101; end
            14'd2767 : begin out <= 64'b0010101100111110001011000001001000100101011010111001110000011011; end
            14'd2768 : begin out <= 64'b1010001110111000001010110000010010101011000011000010101101000010; end
            14'd2769 : begin out <= 64'b0001110000010010000110110011000110101010001010011001010111100011; end
            14'd2770 : begin out <= 64'b1010010111101011001010000000011010100010001001010010101110111001; end
            14'd2771 : begin out <= 64'b0001110010110101101000110011001010100111001011100010101101110000; end
            14'd2772 : begin out <= 64'b1010010100010001001001101100101110101011011110110010101101001111; end
            14'd2773 : begin out <= 64'b0010100101001110101001100100000010101010001100000010000011100001; end
            14'd2774 : begin out <= 64'b0010000001100001101000000010101000100100101100011010100011001100; end
            14'd2775 : begin out <= 64'b1010011001101000101010100000101110100101101101110010100100100111; end
            14'd2776 : begin out <= 64'b0010101001100011000111111111010010101010000010011010100110011110; end
            14'd2777 : begin out <= 64'b0010010110100101001001010111101100101001001000101010010010001111; end
            14'd2778 : begin out <= 64'b1010100101011001001001111101111110100010111011011010001111001110; end
            14'd2779 : begin out <= 64'b0010100111001110001010101101100100101011011111110010101111011111; end
            14'd2780 : begin out <= 64'b0010001000011100101010001111011100101001100111011010101000000101; end
            14'd2781 : begin out <= 64'b1010011101111001101010010111100000100010111111011010100111001101; end
            14'd2782 : begin out <= 64'b0010101000010100101001000101000000010111100100110010100010011100; end
            14'd2783 : begin out <= 64'b0010101101101110101000100011000000101000110011110010101101101010; end
            14'd2784 : begin out <= 64'b1010101011111001101011000011010110011110001101010010100100010000; end
            14'd2785 : begin out <= 64'b1010000000111011100110101011011010101011010110000001101010011011; end
            14'd2786 : begin out <= 64'b1010000010000010101001000101010110100110011100000010010101010010; end
            14'd2787 : begin out <= 64'b0010101010111100101000001010010010100000100010011010011000111011; end
            14'd2788 : begin out <= 64'b1010001110110010001001100110000100101001111010001010001100000111; end
            14'd2789 : begin out <= 64'b1010000111100100101010000001010110100101000101111010100010101000; end
            14'd2790 : begin out <= 64'b1010010010100010001010110101111010100011111000001010101011010000; end
            14'd2791 : begin out <= 64'b1010001101101000101010001100010100101010111001011010101000110101; end
            14'd2792 : begin out <= 64'b0010101101111001001010000110000110101001110000000010000100100101; end
            14'd2793 : begin out <= 64'b0010000001110110101010000111000100101001110100000010011111010000; end
            14'd2794 : begin out <= 64'b0010010001111001001001001000010000101011000110101010011001011011; end
            14'd2795 : begin out <= 64'b1010011100010110001000110110100010101011110000000010101011001100; end
            14'd2796 : begin out <= 64'b0010100111101011101010001001011100101011001100110010001110001001; end
            14'd2797 : begin out <= 64'b1001110010111110001010011100110000101010100111110001100000011011; end
            14'd2798 : begin out <= 64'b0010101010000111101001101101111000101010011101001010011011101110; end
            14'd2799 : begin out <= 64'b1010101011100111001010101010110000101000110110001010011101111100; end
            14'd2800 : begin out <= 64'b1010101110001111001001111010100100101010100001101001111010110100; end
            14'd2801 : begin out <= 64'b0010010011001110001010101101100110100101000100000010011101010110; end
            14'd2802 : begin out <= 64'b1010001000110000101001100101010110011111000001011010100011000011; end
            14'd2803 : begin out <= 64'b0010100111111000001010111101101000100110000100011010100110010001; end
            14'd2804 : begin out <= 64'b1010011001001000001010101100001000101010011011100010100110000000; end
            14'd2805 : begin out <= 64'b0010100101001100100111010000100000101010111011001010010010001011; end
            14'd2806 : begin out <= 64'b1010100010010111100111111100101010100101110101110010100110000111; end
            14'd2807 : begin out <= 64'b1010101111010100101001100011100110101011100110101010100110100101; end
            14'd2808 : begin out <= 64'b0010101000001110001010000011010100101000101010110010011110101111; end
            14'd2809 : begin out <= 64'b1001111100100110001010001010101010100010001110101010101101000010; end
            14'd2810 : begin out <= 64'b0001111010001101101001001001010010100110110100011010010010101001; end
            14'd2811 : begin out <= 64'b0010010100000111001010011101111110101011100011000010000110101100; end
            14'd2812 : begin out <= 64'b0010101010011111001001111010001000011110011000010001111010010011; end
            14'd2813 : begin out <= 64'b1010010001001000001001110010000000100110110110010010101011101000; end
            14'd2814 : begin out <= 64'b1010000111000011101000001010110100101001010000110010101010110000; end
            14'd2815 : begin out <= 64'b1010101000101100101000110101010000101010100010100010101101000000; end
            14'd2816 : begin out <= 64'b0010100010110110101001000101100000101001000100001010101000001110; end
            14'd2817 : begin out <= 64'b1010010000110000101001101101111110100011010001101010101111001100; end
            14'd2818 : begin out <= 64'b1001110000001101001010010010011110100100011101010010101011010001; end
            14'd2819 : begin out <= 64'b0010100001001101001001001011000100100111000111011010100101001101; end
            14'd2820 : begin out <= 64'b1010100100010101000111001110111000011000000001010010010000110111; end
            14'd2821 : begin out <= 64'b1001110000001101001001110001000010101000000011111010101101010101; end
            14'd2822 : begin out <= 64'b1010101101000010100110101111000100100111001001011010100100001110; end
            14'd2823 : begin out <= 64'b0010011101001010101001110110001100101010101010000010010110111111; end
            14'd2824 : begin out <= 64'b0001101010011000001000001100001000101010000110010010011100110010; end
            14'd2825 : begin out <= 64'b1010011100011111101001011011100100101010110011101010100001011101; end
            14'd2826 : begin out <= 64'b0010100110100010001010111111011110101001100001000010100111110000; end
            14'd2827 : begin out <= 64'b1010101000001101101010111001110010101001101011110010100110000001; end
            14'd2828 : begin out <= 64'b1010010000010111001010111001100110100111111001000000100001010110; end
            14'd2829 : begin out <= 64'b0010100001010010001010010010111100011110100010100010101101000100; end
            14'd2830 : begin out <= 64'b1010011101011110001010111110011100101001100001010010101110010110; end
            14'd2831 : begin out <= 64'b1010010001111000101000100111100110011101011111011010101100000010; end
            14'd2832 : begin out <= 64'b0010010100011101101010100110110100101010001101101010101000110010; end
            14'd2833 : begin out <= 64'b1010011111011111101010011111011110101001000111010010100101100110; end
            14'd2834 : begin out <= 64'b1010011011010110101010111011111000100010000010000010101000011000; end
            14'd2835 : begin out <= 64'b0010100010010101101010111010110100100111010001010010011010011011; end
            14'd2836 : begin out <= 64'b1010000001001110101010000010000110100111010001000010010000100101; end
            14'd2837 : begin out <= 64'b1010011000001010000111011010001000101000111000100001111001111000; end
            14'd2838 : begin out <= 64'b1010101110001111101001111111000100100011100110001010010100010111; end
            14'd2839 : begin out <= 64'b1001110000110010101010101001101100011100101000111010010000001111; end
            14'd2840 : begin out <= 64'b1010010110100010101010011000111000100001110100011010101000101101; end
            14'd2841 : begin out <= 64'b1010100100111010000111111100001000101010111001110010100011100101; end
            14'd2842 : begin out <= 64'b0010100100101110001001000100101110100011100111111010101000001101; end
            14'd2843 : begin out <= 64'b1010100001100011001010000101010110100000100001111010100111000000; end
            14'd2844 : begin out <= 64'b0010100101001011000111101001110010101001111001000010010101000100; end
            14'd2845 : begin out <= 64'b1010010111000001101001101100011110100100110001011010101101101101; end
            14'd2846 : begin out <= 64'b0010100010111001101001110010110010100111011001101010001111000100; end
            14'd2847 : begin out <= 64'b1001110101010000100101001001000000101001010001110010100001110001; end
            14'd2848 : begin out <= 64'b0010011110000000101010101110111110101001000100000010100101110100; end
            14'd2849 : begin out <= 64'b1001111000111100101010000100101000100000011101011010100111011011; end
            14'd2850 : begin out <= 64'b1010010101100110001010001000011010100111011111011010100100101111; end
            14'd2851 : begin out <= 64'b1010101011000001000111000000011110101011010101110010110000000110; end
            14'd2852 : begin out <= 64'b1010100000110110101001010001000000101001011000110001101101001100; end
            14'd2853 : begin out <= 64'b1010011110110011101000011110010010011001110100001010011101101001; end
            14'd2854 : begin out <= 64'b0001110110011010101000101111001010101010010110100010100110100010; end
            14'd2855 : begin out <= 64'b1001100101110011101001010011011010101000001100001010100110010001; end
            14'd2856 : begin out <= 64'b0010100110011100001001011110111000101011001110100001101101101100; end
            14'd2857 : begin out <= 64'b0010100101000110101010000011010000101011111011110010011101011111; end
            14'd2858 : begin out <= 64'b0010101101111101001000111101101000011010010001101010101101101100; end
            14'd2859 : begin out <= 64'b0010011011101011101010010110111000101001110101010010100010100101; end
            14'd2860 : begin out <= 64'b1010001111011000001010100110100010101000001000000001100010110011; end
            14'd2861 : begin out <= 64'b0010001110101011100110011110000000101001001110000010100110101000; end
            14'd2862 : begin out <= 64'b1010010001101101101010111111110010100000100101111010101110010011; end
            14'd2863 : begin out <= 64'b1010101000101111001010010001101110100010111011011010101100101011; end
            14'd2864 : begin out <= 64'b1010101000010000001010110010010100100101111101101010101011011000; end
            14'd2865 : begin out <= 64'b0010010001011001001010100101111110100101100011110010001110000011; end
            14'd2866 : begin out <= 64'b0010101110011011101010011111100000101011011000001010101111010001; end
            14'd2867 : begin out <= 64'b0010000100000011101001110011010110100101110000001010100000111101; end
            14'd2868 : begin out <= 64'b1001111010000100001001010001100110100101110010011010011101000010; end
            14'd2869 : begin out <= 64'b0001100010011010101000110010000010101000111111111010101000011100; end
            14'd2870 : begin out <= 64'b0010101001001111101001000011101000100110010011111010100010111000; end
            14'd2871 : begin out <= 64'b0010100101010010001010101010001010101010010110110010001000111011; end
            14'd2872 : begin out <= 64'b1010010111001011000110010110101110101010101100111010100001101110; end
            14'd2873 : begin out <= 64'b0010000011101001000111100110100110101000011110101010101010101100; end
            14'd2874 : begin out <= 64'b0010011000000110101000111011010010101000010111010010100011101110; end
            14'd2875 : begin out <= 64'b1010100001001011001010100010101010100001011011010010100000100100; end
            14'd2876 : begin out <= 64'b0010011111110010000100010000100010101011100011010010010001001100; end
            14'd2877 : begin out <= 64'b0010100101010000101010111101110100011010011100001010010101101101; end
            14'd2878 : begin out <= 64'b0010010010111000001010001001000000101001101100010001101001011101; end
            14'd2879 : begin out <= 64'b0010101101101100101010000110001010101010011000100010001111001101; end
            14'd2880 : begin out <= 64'b0010101110100110001010010110010100011101110010101010100111000010; end
            14'd2881 : begin out <= 64'b1010011000010110001010110110110110101000000111111010100001011110; end
            14'd2882 : begin out <= 64'b0010011011000001001010100000100010101011011011010010010101100110; end
            14'd2883 : begin out <= 64'b1010100011110000001010101011111010100111101110000010101010110001; end
            14'd2884 : begin out <= 64'b0010100000001001101010100000100110100110110111110010001001001111; end
            14'd2885 : begin out <= 64'b0010010111100011101001000010110100100111010010001010001011010000; end
            14'd2886 : begin out <= 64'b1010100101110011101000010011110100101000100101000001101110001110; end
            14'd2887 : begin out <= 64'b1010010010011000101010101001111000100111101011101010100111000010; end
            14'd2888 : begin out <= 64'b0010100000000111101010011101100010100011000001101010010011010100; end
            14'd2889 : begin out <= 64'b0010101110110011001010001001100000101001101011101010010111000101; end
            14'd2890 : begin out <= 64'b0010100011011100101001101000000010100101010011101010100011000110; end
            14'd2891 : begin out <= 64'b1010101001101111101010010000001010001101011101001010101011110100; end
            14'd2892 : begin out <= 64'b0010010011111100101010100011001110100000011011111010101101010000; end
            14'd2893 : begin out <= 64'b0010010100000001101001100101110000101010001101110010101111000111; end
            14'd2894 : begin out <= 64'b1010100111101100101001000101101010100111111010110010101101100000; end
            14'd2895 : begin out <= 64'b0010100111110110001010000101101110101010000100001010011010001111; end
            14'd2896 : begin out <= 64'b0010101100101010101010001101011010100000001001011010101101110001; end
            14'd2897 : begin out <= 64'b0010010011001101101000000101110000100000011001010010011000111011; end
            14'd2898 : begin out <= 64'b0001100100011011001010110101110010100011001111111001100010110101; end
            14'd2899 : begin out <= 64'b0010010010000000001000101010110000100110000100110010010010110111; end
            14'd2900 : begin out <= 64'b0010100101001101101000001101111100101000100100010001111101010111; end
            14'd2901 : begin out <= 64'b0010100011000000101000110010000100101000010010000001110010111101; end
            14'd2902 : begin out <= 64'b0010000001110111000111011011110000101011000111100010100110010000; end
            14'd2903 : begin out <= 64'b0010011000001010101010010101011110101000001010100010011110001011; end
            14'd2904 : begin out <= 64'b0010100111111100100110110111010100101010101011100010101111110110; end
            14'd2905 : begin out <= 64'b1010000001011100101000100100100110101001000011000010011010111111; end
            14'd2906 : begin out <= 64'b0010101001011010001010011000000100101010000001100010010000101101; end
            14'd2907 : begin out <= 64'b0010000010010101001010110000000110101011001010001010001111100000; end
            14'd2908 : begin out <= 64'b0001110110100001001010011000010110101000111100000010101111011001; end
            14'd2909 : begin out <= 64'b1010101000000100001001010101101000011101000000001010100101011000; end
            14'd2910 : begin out <= 64'b0010010000101111101010100100011110101011010101111010101000010110; end
            14'd2911 : begin out <= 64'b0001110001100100001010010001110110101001110111000010101011101000; end
            14'd2912 : begin out <= 64'b0001100110010100001010011011101010100110101100010010101111011000; end
            14'd2913 : begin out <= 64'b1010100101011001101001001111010100101011101001000001001100100010; end
            14'd2914 : begin out <= 64'b0010011111001100101010000101001010101010100101101010100111110110; end
            14'd2915 : begin out <= 64'b0010100101000110000111000111001100101011111111110010000010001111; end
            14'd2916 : begin out <= 64'b1001110000001101001010011100011010100000001011110010011011111100; end
            14'd2917 : begin out <= 64'b0010001010010110101000100001101000101001110000101010010100111111; end
            14'd2918 : begin out <= 64'b1010010111000110000111001101011100100001000100000010010001000100; end
            14'd2919 : begin out <= 64'b0010101011010000100111010011100110100000010110100001011110111101; end
            14'd2920 : begin out <= 64'b1001011110010001101010011101110110101000011100101010101001110100; end
            14'd2921 : begin out <= 64'b0010100010100010000110010010100010101000101101101010100000110110; end
            14'd2922 : begin out <= 64'b1010011100001101001001101110110010100110111010101010010000011110; end
            14'd2923 : begin out <= 64'b1010101000000100001001001001111000010010010101110010010001000100; end
            14'd2924 : begin out <= 64'b1000111000000001101010011111011000100000111000101010010110000110; end
            14'd2925 : begin out <= 64'b0010010110001010001001010011011000101010001111000010100111001111; end
            14'd2926 : begin out <= 64'b1010101011100110100110010111111000100001011001010001111110010001; end
            14'd2927 : begin out <= 64'b1010100000000111001001111000001110101000111101011010100011101111; end
            14'd2928 : begin out <= 64'b0010101101010000000110111000111110101011111111000010100110100011; end
            14'd2929 : begin out <= 64'b0010101010111100001001100011110110101010001100011010001010110010; end
            14'd2930 : begin out <= 64'b1010010110111000001010000000100100100111101011011010100101001111; end
            14'd2931 : begin out <= 64'b1010100001000001101010001111101100100101111101111010100101111010; end
            14'd2932 : begin out <= 64'b0010100001101110001001000011011010101001111011001001011111100000; end
            14'd2933 : begin out <= 64'b0010011111010100101010001011111110101010100010101010000110110111; end
            14'd2934 : begin out <= 64'b0010101100100100001001000011101000101011110011101010100100101011; end
            14'd2935 : begin out <= 64'b0010010101111010001010111000101000101000110011110010101000111100; end
            14'd2936 : begin out <= 64'b0001110101001001101000100010110100011101111110101010000010110010; end
            14'd2937 : begin out <= 64'b0010011001111110100010000001000110100111111110001010011010110010; end
            14'd2938 : begin out <= 64'b0010100111100000101000011111010010101000010000001010100011101111; end
            14'd2939 : begin out <= 64'b1010011101111000101000011100010010011111001010100010100010111100; end
            14'd2940 : begin out <= 64'b0010100111011010001010101010100110100110011000111010011100001100; end
            14'd2941 : begin out <= 64'b0010100110011010101001111100100010100100001111110010101010111101; end
            14'd2942 : begin out <= 64'b1010011010111000101001111000100110101011000000010010001010001111; end
            14'd2943 : begin out <= 64'b1010100111101001101000100000011110100111111010110001110001100010; end
            14'd2944 : begin out <= 64'b1010101000000111101001100010001010100000101011000010101011101100; end
            14'd2945 : begin out <= 64'b0010101000101110001001111010010010101011110001111010011011100111; end
            14'd2946 : begin out <= 64'b1010000101111101101010001101000010101000001100011010100011101110; end
            14'd2947 : begin out <= 64'b0001101010001001101001110001010100101000101111000010101011110011; end
            14'd2948 : begin out <= 64'b1001110110000110101001101001110110011100100011111010001100111100; end
            14'd2949 : begin out <= 64'b1010010110101101101001010000100100101000000010001010011001001100; end
            14'd2950 : begin out <= 64'b0010100011010100101001101101100010100101100101011001111100100111; end
            14'd2951 : begin out <= 64'b1010010000111111101001111010110010101000010100111010000100110100; end
            14'd2952 : begin out <= 64'b1001101000001011101010101000100000101010011111010010011000110100; end
            14'd2953 : begin out <= 64'b0010010111110101100010010001010100101011000001100001000010100000; end
            14'd2954 : begin out <= 64'b0010101011000001101001111101011010101000010110010010010100000010; end
            14'd2955 : begin out <= 64'b1010010010010110001001001011100100010011100101001001110100011111; end
            14'd2956 : begin out <= 64'b1010010101110010001010110010110110101000001010011010011111110100; end
            14'd2957 : begin out <= 64'b1010101110110011101010111101101100101001000010000001111110000110; end
            14'd2958 : begin out <= 64'b1010101101001001001000001110011110101000010001010010010010010110; end
            14'd2959 : begin out <= 64'b0010100000000010001010100100001110101010000010001010100101111000; end
            14'd2960 : begin out <= 64'b1010011000110110101010010001001100101010000101011010001010110001; end
            14'd2961 : begin out <= 64'b0010011111101010101010001010010100100111011001010010101001011100; end
            14'd2962 : begin out <= 64'b1010101111001010001010000110110000100010101100110010010101001111; end
            14'd2963 : begin out <= 64'b0010101101011101101010101111011100011111101111100010010011110001; end
            14'd2964 : begin out <= 64'b0010100110000001101000011100010100100111111011101010100101000011; end
            14'd2965 : begin out <= 64'b1010100000000101001001000111000110011011110110011010010010001000; end
            14'd2966 : begin out <= 64'b0010010111101100001001001001100100101010010011001010011010110000; end
            14'd2967 : begin out <= 64'b1010100001110110001000111001011010101011010000011010100100000001; end
            14'd2968 : begin out <= 64'b0010011001110000101010000100000110101010100011111010100111011010; end
            14'd2969 : begin out <= 64'b1010011111110011101010110101001110101001101011011010100100100011; end
            14'd2970 : begin out <= 64'b1010010000011010101010001001100110101010100001111010010010110001; end
            14'd2971 : begin out <= 64'b0010010001010010000110011101110010101001101000000010100000010001; end
            14'd2972 : begin out <= 64'b0010100001000101101010100001011110100111100101000001010101100111; end
            14'd2973 : begin out <= 64'b0010000010100001001000110010100000101000101111001010001110001000; end
            14'd2974 : begin out <= 64'b1010100101111011001001111010101010100000111110100010000110010101; end
            14'd2975 : begin out <= 64'b1010010110001100101010101110110110101000000100111010100000100100; end
            14'd2976 : begin out <= 64'b1010001101110111001000100101100100100011001111101010011111110100; end
            14'd2977 : begin out <= 64'b0010100010101110001001010011111010101010110110000010101010010110; end
            14'd2978 : begin out <= 64'b0010101101010000101010111110101110100110100101111010100100111001; end
            14'd2979 : begin out <= 64'b0001010100010001101010000110110100100101110101100010011001100111; end
            14'd2980 : begin out <= 64'b0010001101011001001010001010100010101011001001111010010111010011; end
            14'd2981 : begin out <= 64'b0010011100011101101000111000111010101010110001001010010010111000; end
            14'd2982 : begin out <= 64'b1001100111010011101001000100111100101010000111110010011101001111; end
            14'd2983 : begin out <= 64'b0010101001101111101001001101101110100111101000110010010010000101; end
            14'd2984 : begin out <= 64'b1010101010000001001010110100000010101010000001000010100101101001; end
            14'd2985 : begin out <= 64'b0010010111010111100101011101110000100101100000011010010011110010; end
            14'd2986 : begin out <= 64'b0001111001001011101001111100011100011011100110101010101111010110; end
            14'd2987 : begin out <= 64'b0010100000011111101010011111100110101000111010100010010011000111; end
            14'd2988 : begin out <= 64'b1010101111010010001001111101101110101000011010101001111000111111; end
            14'd2989 : begin out <= 64'b0010100011001010001001111110111100011000011000010010101110110010; end
            14'd2990 : begin out <= 64'b1010100001101000001000111000011010011100101000100010100010001100; end
            14'd2991 : begin out <= 64'b0010100011101000000111111000010010011010100011100010101011100110; end
            14'd2992 : begin out <= 64'b1010000001000101101010010000110100101011101010100001110110010110; end
            14'd2993 : begin out <= 64'b1010001011111011101010100010110010100010011001110010000101011101; end
            14'd2994 : begin out <= 64'b0001010000110010101010110111001010101000101010000010101100010110; end
            14'd2995 : begin out <= 64'b1010011101011010101010100001011100101000011101101010000000010100; end
            14'd2996 : begin out <= 64'b0010011100000000001001110101101100101010111101101010010001000101; end
            14'd2997 : begin out <= 64'b0010100010101111001010110011110110100100011000010010101001111001; end
            14'd2998 : begin out <= 64'b1010011111011110100100011101010110101000001111111010100100100010; end
            14'd2999 : begin out <= 64'b1000001111010010001010010010001000101000011101110010100010000001; end
            14'd3000 : begin out <= 64'b0010100101111011101001111110100110100000101110000001111111000001; end
            14'd3001 : begin out <= 64'b1001101000010001101010000010000110101010111001111010101000110011; end
            14'd3002 : begin out <= 64'b0010101001001101100110110010001000100111100101111010100011111000; end
            14'd3003 : begin out <= 64'b0010011011101100000110001001000000101010001000101010101001101101; end
            14'd3004 : begin out <= 64'b0010011001011111001001100101010000101011111100110001110000011101; end
            14'd3005 : begin out <= 64'b1001010111001111000111000010110100101011011110010010101011000000; end
            14'd3006 : begin out <= 64'b0010100000111100001001001010100000100011110011110001010100110000; end
            14'd3007 : begin out <= 64'b0010010000010001000110110111001000101010010001111010000010100000; end
            14'd3008 : begin out <= 64'b0010100011111000101001111010001010101010111011100010001010001111; end
            14'd3009 : begin out <= 64'b1010101100101010101001111101001010101010000110010010100000100100; end
            14'd3010 : begin out <= 64'b1010000011101100001010111111011000101001010010001010100000011111; end
            14'd3011 : begin out <= 64'b0010101110011110100011100110001010100100111110010010101000101001; end
            14'd3012 : begin out <= 64'b1010001101101011001001000101110000101011011000101010100100100101; end
            14'd3013 : begin out <= 64'b1010101001001001001010110010101010101011111100101010100011011011; end
            14'd3014 : begin out <= 64'b0010100010000000100111001110110010100010111011110001110011001010; end
            14'd3015 : begin out <= 64'b1001110010110101001010100011000100100100011110101000100000110111; end
            14'd3016 : begin out <= 64'b0010101100000000001001011100011000011111000001010010010111010101; end
            14'd3017 : begin out <= 64'b1010101101011111000110011010110000101011111110000001110001101001; end
            14'd3018 : begin out <= 64'b1010101100000111001001111101100110010100000001111010101011101001; end
            14'd3019 : begin out <= 64'b0010011100101110101010100111110100101010011110010010000100010001; end
            14'd3020 : begin out <= 64'b1010101100000111001000011100010000011010101110001010011110001110; end
            14'd3021 : begin out <= 64'b1001011011010000001010110000001000100100100101111010101001101100; end
            14'd3022 : begin out <= 64'b0010010110000110000111110111111010101001100011110010101111100100; end
            14'd3023 : begin out <= 64'b1010001101001101101010001100011010101000001100001010010110011100; end
            14'd3024 : begin out <= 64'b0010011110111000101010011000110110100100011100110010100011001001; end
            14'd3025 : begin out <= 64'b0010000110011110001010001100011100010100100101010010101100110001; end
            14'd3026 : begin out <= 64'b0010010001010011101010100001111010100111011011110010011100100000; end
            14'd3027 : begin out <= 64'b0010000000111001001010101010010000011100111101010010100010110000; end
            14'd3028 : begin out <= 64'b0010010111011101001001101110011110101000010101100010011001001011; end
            14'd3029 : begin out <= 64'b1010010101100110101000000000000110101000111001000010110000001111; end
            14'd3030 : begin out <= 64'b0010000011001001001000110101011010100100010010001010101010111011; end
            14'd3031 : begin out <= 64'b0010010011111100001001010111110110100100101101101010100101101100; end
            14'd3032 : begin out <= 64'b0010001010111000101010011011101110101001011100101010001111111100; end
            14'd3033 : begin out <= 64'b0010100010101011100111100100110100101010011000111001011111100111; end
            14'd3034 : begin out <= 64'b1001101110000101101000100101010000010001010011100010100100010111; end
            14'd3035 : begin out <= 64'b0010010111010101001010010111101010100111110101000010100000111001; end
            14'd3036 : begin out <= 64'b0010101011111000101010111111110010100111010110011010011001011100; end
            14'd3037 : begin out <= 64'b1010100010110110100111100001110000101011111010011010110000001000; end
            14'd3038 : begin out <= 64'b1010101101100111001010110011100100100110100111011010101000111011; end
            14'd3039 : begin out <= 64'b1010101010111101101010010100110010101010100110110010101101001110; end
            14'd3040 : begin out <= 64'b0010100100111111001010100110110110100110001011110010010101100111; end
            14'd3041 : begin out <= 64'b1010101001110101101001101011000000100001110100111010100000110011; end
            14'd3042 : begin out <= 64'b1001111011011010001010111001111110101011011100111010100101101011; end
            14'd3043 : begin out <= 64'b0010001100101010100110011011100100101000111101010010001011100001; end
            14'd3044 : begin out <= 64'b0010001111001011001010101101001010101001010010000010010000100101; end
            14'd3045 : begin out <= 64'b1010101011011000001010100000111010011001100010011010000001000011; end
            14'd3046 : begin out <= 64'b0010000111010101001010010010110100100110000011100010100011010110; end
            14'd3047 : begin out <= 64'b0010101111101001101000100110000100100101001101110010100110110001; end
            14'd3048 : begin out <= 64'b0010100011001101101010101000100100101000110110000010101101000110; end
            14'd3049 : begin out <= 64'b0001111110000000101010110001001110101000010100001010101011110111; end
            14'd3050 : begin out <= 64'b0010101000010111001000010111100100100111100111111001101100000100; end
            14'd3051 : begin out <= 64'b0010100010000011001000111000010010100101010101000010011011000101; end
            14'd3052 : begin out <= 64'b1010100011101110101010111100011100101000111011101010011010001011; end
            14'd3053 : begin out <= 64'b1001110111010110001001011110011010101000111100010010100111101101; end
            14'd3054 : begin out <= 64'b0010100001111110001010111011110010100100010010010010011011010100; end
            14'd3055 : begin out <= 64'b1001111001100000101000000111000000011111000100011010100111111011; end
            14'd3056 : begin out <= 64'b1010100000110000000110111100001000101011101110010010011111101111; end
            14'd3057 : begin out <= 64'b0001001110111000001010000100110010100011000101011010101000101101; end
            14'd3058 : begin out <= 64'b1010101000000111001000110011100010101000100011001010011100100001; end
            14'd3059 : begin out <= 64'b0010101110100110101010000100011010101001110111111010101000111000; end
            14'd3060 : begin out <= 64'b0010100101111101001000100111110100101000100100000010000011110100; end
            14'd3061 : begin out <= 64'b0001111001101001001001101011101000100111001110011010101001001010; end
            14'd3062 : begin out <= 64'b1010010100100110001010001111001100100110011110100010011111000011; end
            14'd3063 : begin out <= 64'b0010011111001011001010110000001100011000000001110010100100101010; end
            14'd3064 : begin out <= 64'b0010100111001011001010110000000100011111100001100010010100010001; end
            14'd3065 : begin out <= 64'b1010010011001100101010000000111010101000011111000010100000100000; end
            14'd3066 : begin out <= 64'b1010011100101000100110000010100010101011100000110010110000000110; end
            14'd3067 : begin out <= 64'b1010101110010111001000011110011110101001000100110010101010100111; end
            14'd3068 : begin out <= 64'b0010101000011011101010000111011110011011010001010010010111001010; end
            14'd3069 : begin out <= 64'b1001111011001001101001111101000000101001001001101010001000000101; end
            14'd3070 : begin out <= 64'b1010010111001111101010010101110100100100010111000010101010110000; end
            14'd3071 : begin out <= 64'b1001111000001011101010100001000010101001101100111010010101010010; end
            14'd3072 : begin out <= 64'b1010000110101001001010111101010000101010010101110010011001101100; end
            14'd3073 : begin out <= 64'b1010100101000111101010110101001010101001010010101010100010000010; end
            14'd3074 : begin out <= 64'b0001011111001011101001110110000000011100111010000010101011000001; end
            14'd3075 : begin out <= 64'b1010100000011010001010111110111000100001001011000010100100111110; end
            14'd3076 : begin out <= 64'b1010010010100110101000011111001110100010111110001010100110110100; end
            14'd3077 : begin out <= 64'b1010001111110101001001011001011010100101001100010010101101101000; end
            14'd3078 : begin out <= 64'b1010101010011000001010011101101110101001110101010001110010111111; end
            14'd3079 : begin out <= 64'b0010100010100111001010101100111100101001101111110010101101101110; end
            14'd3080 : begin out <= 64'b0010101100111001001010001110001110101010010001110010101100011010; end
            14'd3081 : begin out <= 64'b0010011001000110101001111011100100101010010100000010101101110000; end
            14'd3082 : begin out <= 64'b0010010001010010101010011010110010100011110011000010100111011001; end
            14'd3083 : begin out <= 64'b1010100111100010001001010100111100101011010010001010011011100101; end
            14'd3084 : begin out <= 64'b0010101111001010001010011011100100100100000110100010101000001110; end
            14'd3085 : begin out <= 64'b1010011101100000101001010000111010011111110010101010100110010011; end
            14'd3086 : begin out <= 64'b1010010100101111001000111000001010100010100010110010100000000011; end
            14'd3087 : begin out <= 64'b1010010100101011101001010010100110101001010001011010100010101110; end
            14'd3088 : begin out <= 64'b1010101100110001100101001001110100100111100001010010010111110011; end
            14'd3089 : begin out <= 64'b0010011111010100001010010001110110101000000100101010101100110111; end
            14'd3090 : begin out <= 64'b1010010111110011101010001111000100100110110000010010010111001111; end
            14'd3091 : begin out <= 64'b0001001001000111101010000011001000101010101111001010011100110000; end
            14'd3092 : begin out <= 64'b0010100101100010001010011011000010101000100100100010100100011011; end
            14'd3093 : begin out <= 64'b1001111010111111100111010100100000101011010011100010101001011011; end
            14'd3094 : begin out <= 64'b0010101110011100101010000000100110101011001100011010101100011101; end
            14'd3095 : begin out <= 64'b0010100011111111101001010101000010011000111101001001111110101100; end
            14'd3096 : begin out <= 64'b1010011011010101100001110011100010101010001010011010010110111011; end
            14'd3097 : begin out <= 64'b1010101110011101001010100101000010010110111000000010101101101111; end
            14'd3098 : begin out <= 64'b0010001111000101101000100000101110101001101010100010100111100011; end
            14'd3099 : begin out <= 64'b1010011001010111101010001010000000011010010011011010011001111001; end
            14'd3100 : begin out <= 64'b1010100001100000101010010111110000101010100011001001111001101110; end
            14'd3101 : begin out <= 64'b0001000011010110101010000011110100011100011011001010101100101111; end
            14'd3102 : begin out <= 64'b1010101100011010101000100111011010100001101110010010100010000011; end
            14'd3103 : begin out <= 64'b1010011100101110001010111011110010101011101101101010011100000001; end
            14'd3104 : begin out <= 64'b0010101110110110101010011011001010100110111010101010100110000111; end
            14'd3105 : begin out <= 64'b1001101001111110001000110010001110101000011001001010100010111000; end
            14'd3106 : begin out <= 64'b1010100101100110001000100010111000011100111001000010011001100100; end
            14'd3107 : begin out <= 64'b0010101110011111001001100111110100101001111010110010000001011100; end
            14'd3108 : begin out <= 64'b1010011111001000001001000001010110100001101101110010010101100101; end
            14'd3109 : begin out <= 64'b0010100010000010100111100011101000101010011111000001111110110000; end
            14'd3110 : begin out <= 64'b0010100010001100001010101100100000101001010000111010110000010101; end
            14'd3111 : begin out <= 64'b1010101001011001101010100110101110101011000001011010100001111100; end
            14'd3112 : begin out <= 64'b1010010011011110100101000111010100101011011011010010101100010111; end
            14'd3113 : begin out <= 64'b1010000010001001001010110101001010100111011011101001000010000100; end
            14'd3114 : begin out <= 64'b0010101011111110001001100110011100101010111110100010101000110001; end
            14'd3115 : begin out <= 64'b1010000111110001101001111011001010011101011110111010010010110000; end
            14'd3116 : begin out <= 64'b1010100111101100101010111000101010100110001011001010010010110001; end
            14'd3117 : begin out <= 64'b0010010011001010001001111010101100100111101001100001110100000101; end
            14'd3118 : begin out <= 64'b1010010111110100101001000011100110101011001000111010001111000010; end
            14'd3119 : begin out <= 64'b1010101000111001000111101110011000101001101100101010000111111110; end
            14'd3120 : begin out <= 64'b0010011111011011101001010001100110101100000100100010101100110001; end
            14'd3121 : begin out <= 64'b1010101100001001101000011100011010101001010100111010101011000011; end
            14'd3122 : begin out <= 64'b1010011100101011101010100111101110100001001111011010000110001101; end
            14'd3123 : begin out <= 64'b1010001100001111100111000010100010101011100110010010000001010000; end
            14'd3124 : begin out <= 64'b0010011000110111001000100110111100100111010110011010110000000000; end
            14'd3125 : begin out <= 64'b1010101000010110001000100101011010101001111001101010101001000111; end
            14'd3126 : begin out <= 64'b0010000111000011001010001011101000101001100010001010101000011000; end
            14'd3127 : begin out <= 64'b1010101110011100001001101001011100101011010001101010101000100101; end
            14'd3128 : begin out <= 64'b0010000100011011101001001010100110101001100011010010011100101001; end
            14'd3129 : begin out <= 64'b1010100000111000001010010011101100001111001111101010001000011100; end
            14'd3130 : begin out <= 64'b0010101111001100001001111001110100101001101001011010011011000000; end
            14'd3131 : begin out <= 64'b1010010011100011000110000100001100100111010110000010011111011010; end
            14'd3132 : begin out <= 64'b1010101100001001001001100100011110101001101101100010000101001011; end
            14'd3133 : begin out <= 64'b0010101110111100001010001101011100100011000011100010000011000100; end
            14'd3134 : begin out <= 64'b1010010110100000101010011101000100101011001001100010101000100001; end
            14'd3135 : begin out <= 64'b0010011001101011001010001100010100010100001011111010001100101111; end
            14'd3136 : begin out <= 64'b1010101001101001101010001000000110011100101100000010011100001110; end
            14'd3137 : begin out <= 64'b0010011110000011001010101111010000101000101001101001001011110100; end
            14'd3138 : begin out <= 64'b0001010000111011101010000001001010100011110011000010010011011111; end
            14'd3139 : begin out <= 64'b0010101000100101001010011011000000101000000000100010011010011010; end
            14'd3140 : begin out <= 64'b1010100011001100101001101111101000101010110101110001111100011010; end
            14'd3141 : begin out <= 64'b1010010001101001001010000011001110100110000000101010100011110110; end
            14'd3142 : begin out <= 64'b1010101001000101101000011101110110101001001010010010100100000010; end
            14'd3143 : begin out <= 64'b0010011010011110001000001101111100100100000100110010000001000111; end
            14'd3144 : begin out <= 64'b0010001001111101101010001001011100101001111110101010000111100111; end
            14'd3145 : begin out <= 64'b1001101010001101001010010100010110011000110011001010101111000011; end
            14'd3146 : begin out <= 64'b0010101110101100101001010001000110100001001010010010000100111101; end
            14'd3147 : begin out <= 64'b0010010011001101001010000011100010101100000000011001110011010111; end
            14'd3148 : begin out <= 64'b0010000111111100101000100110110010100110000101000010011001001101; end
            14'd3149 : begin out <= 64'b0010011100100111100111011100101000101010011010111010101000000110; end
            14'd3150 : begin out <= 64'b1010101110100001101000111011101000100101100000101010011011111110; end
            14'd3151 : begin out <= 64'b0010011000110011101010101100010100100110111111100010100110110101; end
            14'd3152 : begin out <= 64'b1010000010011101001010001011000010101010010010011001110111110111; end
            14'd3153 : begin out <= 64'b0010100110001001101010110000011000101010010100011010100111011001; end
            14'd3154 : begin out <= 64'b1010010001001011000111111101110100101011010001101010101011110011; end
            14'd3155 : begin out <= 64'b0010100110011111101001100001101110011110010111101010100101001011; end
            14'd3156 : begin out <= 64'b1010010111110001101010010110111100101010101001010010010111010001; end
            14'd3157 : begin out <= 64'b1010101010010111000101110001101110100011011111100010101111000010; end
            14'd3158 : begin out <= 64'b1010100010001011101000100001111000100010010101011010101000000010; end
            14'd3159 : begin out <= 64'b0010010010011110100110001111011010101010000011110010101000100000; end
            14'd3160 : begin out <= 64'b1010101100110101101000110101110100011010010100100010100100011100; end
            14'd3161 : begin out <= 64'b0010010111011000001000011101001110101011111000110010100111001011; end
            14'd3162 : begin out <= 64'b1010000000101101101010011100011110100110100011010010011101101001; end
            14'd3163 : begin out <= 64'b0010100100100000101001000101110010100111001101010010000011011010; end
            14'd3164 : begin out <= 64'b0010100010001000001011000000000010100000100001111010000001100100; end
            14'd3165 : begin out <= 64'b0010010110101000101010101111111110101000010010010010000011000100; end
            14'd3166 : begin out <= 64'b1010011110011100001001000000000110100110000010100010101111110001; end
            14'd3167 : begin out <= 64'b0010001011000100101010110001011100101011100111110010100101011010; end
            14'd3168 : begin out <= 64'b1010101011010000101000111110001100101011000111101010001011100101; end
            14'd3169 : begin out <= 64'b0010100010100001101000011111110100100100111001101010100001011010; end
            14'd3170 : begin out <= 64'b1010101101000010001010111011011100101000111101011010101111101011; end
            14'd3171 : begin out <= 64'b1010101111010011001010110001000110101000000101100001111110000110; end
            14'd3172 : begin out <= 64'b0010101100101001000110001000011000100111000000001001110110010000; end
            14'd3173 : begin out <= 64'b1010011110111110101001110000011000100010001101010010010010001011; end
            14'd3174 : begin out <= 64'b1010001111110101100110001010111100100100100100000010101001101111; end
            14'd3175 : begin out <= 64'b0010000111100110001001011011011100100101000011010010100000101011; end
            14'd3176 : begin out <= 64'b0010000100101100101010101001011010011010000000011010101011010111; end
            14'd3177 : begin out <= 64'b0010101010100001001010100101111010100111000111000001101010100100; end
            14'd3178 : begin out <= 64'b1010100101011011001000110010001110101001000100010010100110110010; end
            14'd3179 : begin out <= 64'b1010100100011101001010101011110110100001100101011010101110011100; end
            14'd3180 : begin out <= 64'b1001111100011010001010011010011000101010011011011010100101101001; end
            14'd3181 : begin out <= 64'b1010011110001011001010111010000100011010110011010010101100010110; end
            14'd3182 : begin out <= 64'b1010010011000110101000100100111110010001110110010010000001111010; end
            14'd3183 : begin out <= 64'b1001111101101110001010011001110100101010011100000010100011101011; end
            14'd3184 : begin out <= 64'b0010011011001011100001011011011110100101101110011010101010110101; end
            14'd3185 : begin out <= 64'b1010101000001101001010100111011000100111010101010010101010001111; end
            14'd3186 : begin out <= 64'b1010010100001100001010111110000010101010001111010010101111000001; end
            14'd3187 : begin out <= 64'b0010010111011010001000111100111000100010001100110010101000111011; end
            14'd3188 : begin out <= 64'b0010100111001000001010110110110010101000111011101010100001101011; end
            14'd3189 : begin out <= 64'b0010101101111000001000010101000000101000101101101010101000101011; end
            14'd3190 : begin out <= 64'b1010011110110101001001010000000100100110010001001010010010001011; end
            14'd3191 : begin out <= 64'b1001110101111111001010010001010010101000011100110010110001000100; end
            14'd3192 : begin out <= 64'b1010101111000110101001101100110100101010100111111001100110101110; end
            14'd3193 : begin out <= 64'b0010011011101100001010000110000000101000000001111010010111100000; end
            14'd3194 : begin out <= 64'b0010101101110010000111011111101100101001100111000010000000010111; end
            14'd3195 : begin out <= 64'b1010101111000110001010110001110000101000011100001010100101110010; end
            14'd3196 : begin out <= 64'b0010101111010010101010000100110000100100001111111010011101011010; end
            14'd3197 : begin out <= 64'b0010001011010001001010100000111010100111101001000010100010001101; end
            14'd3198 : begin out <= 64'b1010010010000110101010110001110010100110110101001010101010110110; end
            14'd3199 : begin out <= 64'b1010010001110000001000101010100010101000101011001010000100101010; end
            14'd3200 : begin out <= 64'b0010010011010111101000010010101000101000000000110010011001001110; end
            14'd3201 : begin out <= 64'b1010011101001101101010011110010110101010100010100010101001110010; end
            14'd3202 : begin out <= 64'b1010100000000110101001100101111010101100001000011010100110000011; end
            14'd3203 : begin out <= 64'b0001101010011010001001110101101110100101011100000010110000010000; end
            14'd3204 : begin out <= 64'b0010010110101010101010011011010110101000001100100010101110100010; end
            14'd3205 : begin out <= 64'b0010101101101010001010111010110100100111010011000010011011011011; end
            14'd3206 : begin out <= 64'b0010101110001100101000011100100100101100000000101010101000001000; end
            14'd3207 : begin out <= 64'b0010100011000001001001010011011110100100001111000010100001000100; end
            14'd3208 : begin out <= 64'b1010101001011000101001010101000000100011110101101010011101000001; end
            14'd3209 : begin out <= 64'b1010011111111100101001110110110110101001001111011010001000110110; end
            14'd3210 : begin out <= 64'b0010100101111011000111011101100110100101111111101010010110110001; end
            14'd3211 : begin out <= 64'b1010101101110100001010010001110010100001011100000010011010001001; end
            14'd3212 : begin out <= 64'b0010100001101011100100111001010110100001110000111001100101001011; end
            14'd3213 : begin out <= 64'b0010010011100111101010110011010000101001000010101010101111011110; end
            14'd3214 : begin out <= 64'b1010100110010001101001111011110110101011001001001010101011100101; end
            14'd3215 : begin out <= 64'b1010001001110110001010100010010110101011110001000010000101000100; end
            14'd3216 : begin out <= 64'b1010001011101110101001001001110010101010001110100010100110000011; end
            14'd3217 : begin out <= 64'b1010010111010111001010000011011000100000111110001010100100110111; end
            14'd3218 : begin out <= 64'b0000111001110001001010110010011010101011101111010010101100001101; end
            14'd3219 : begin out <= 64'b0010011111010111101010011000011110101010111111000010100001010011; end
            14'd3220 : begin out <= 64'b0010001111101011000110010011110110011111111011010001110000100100; end
            14'd3221 : begin out <= 64'b0010010011110011000111001011000000101010110111110010100111100101; end
            14'd3222 : begin out <= 64'b0010101010100001101010101000100010100011010000001010001101000010; end
            14'd3223 : begin out <= 64'b1001000101111100100110101011111110101001010011111010000010100000; end
            14'd3224 : begin out <= 64'b0010001000100101101001101011101010100110110110011010000110111001; end
            14'd3225 : begin out <= 64'b0010101000010000101001110110101000100111100101101001100111101001; end
            14'd3226 : begin out <= 64'b1010000100011011001001001000001100100000000110101010011001001110; end
            14'd3227 : begin out <= 64'b1010100101011011101010000010100010100110010110111001111011010101; end
            14'd3228 : begin out <= 64'b0010100011111000101010101000110000101000101010010010010110000000; end
            14'd3229 : begin out <= 64'b1010010111100111001001011101011010101001110110100010100011111001; end
            14'd3230 : begin out <= 64'b0010011100111010101001010101001010101010100001001010011110111101; end
            14'd3231 : begin out <= 64'b0010101100110111001010000111001100011110101000000010101000101110; end
            14'd3232 : begin out <= 64'b0010100010011011001000011010001110101010100100100010011001110111; end
            14'd3233 : begin out <= 64'b1010001000110010101001010100111100101011100011101010101000100101; end
            14'd3234 : begin out <= 64'b1010100101001111001001001101101100101010010001111010011010111010; end
            14'd3235 : begin out <= 64'b0010100011000110000111100011001000100010111110010010100000000010; end
            14'd3236 : begin out <= 64'b0010100010100110101010110010101110011100111101101010100100101010; end
            14'd3237 : begin out <= 64'b1010100001100110001001010001101010100000111001001010000111000011; end
            14'd3238 : begin out <= 64'b0001110000111100101001111100001100100110101110001010011111001000; end
            14'd3239 : begin out <= 64'b0010100011010000001000000100100010101000001111100010101001011001; end
            14'd3240 : begin out <= 64'b0010100010000010101010111001011010100000001101001010011011101000; end
            14'd3241 : begin out <= 64'b1010011000111101001001001101100000101001100010100010101011101010; end
            14'd3242 : begin out <= 64'b0001011010110000101010000000100010100000101100101010100110000000; end
            14'd3243 : begin out <= 64'b1010010100100000101010111000110110010100011001010010101010001100; end
            14'd3244 : begin out <= 64'b0010010100000000101010110101110100101010110010000001111011101000; end
            14'd3245 : begin out <= 64'b0010101001110000101010000100101110100111100110111010000000110111; end
            14'd3246 : begin out <= 64'b0010101101101011101001101110101100100001111111101010101000110000; end
            14'd3247 : begin out <= 64'b0010101101001000001010001100111100101010110111110010101110000001; end
            14'd3248 : begin out <= 64'b1010100000000110000111110110100000100110000100101010101000111111; end
            14'd3249 : begin out <= 64'b1010101000111001101000101001011010101010010111010010101110100100; end
            14'd3250 : begin out <= 64'b1010100011100110001000011010101000101001010010100010100111111010; end
            14'd3251 : begin out <= 64'b0001110011000010101010001100110110100101110110101010101111111111; end
            14'd3252 : begin out <= 64'b1010100000101101001001100100000110100111010011111010101011010000; end
            14'd3253 : begin out <= 64'b0001111101110010101010000110011000101010010110010010011111100010; end
            14'd3254 : begin out <= 64'b1010100001011011101001011100101010101010001011011010010100110110; end
            14'd3255 : begin out <= 64'b1010100010100000001010100110101000101001000000000010101111010000; end
            14'd3256 : begin out <= 64'b1010100011001101101001000001110000100100010101011010011101110000; end
            14'd3257 : begin out <= 64'b1010010000001110101010010110110010100110001001010010010000101001; end
            14'd3258 : begin out <= 64'b1010101011101100001010001101001000101000111100111010100110100110; end
            14'd3259 : begin out <= 64'b0010100000001101001001101010010000100101111011010001011000100011; end
            14'd3260 : begin out <= 64'b0010100001001101001000110100110100101000001011111010100110011110; end
            14'd3261 : begin out <= 64'b1001111111010100000111011011101010101000110011011010010010001010; end
            14'd3262 : begin out <= 64'b0010011101010010101001110101110110101000000010111010100001001011; end
            14'd3263 : begin out <= 64'b1010010011110000001001011111111100100010100110110010101101010101; end
            14'd3264 : begin out <= 64'b1010101101001010001001010010000110011011110010111010001001100100; end
            14'd3265 : begin out <= 64'b1010100000000001101001001000000000011101000000100010010101011100; end
            14'd3266 : begin out <= 64'b1010101101100101001001100000101000101001000110101010100111011000; end
            14'd3267 : begin out <= 64'b1010101010110100101010011001111000100100111111000010100100010101; end
            14'd3268 : begin out <= 64'b1010100101001110100111010110111000101000001110010010010111000001; end
            14'd3269 : begin out <= 64'b1010011111100011001010010111011000101010101000000010101001111100; end
            14'd3270 : begin out <= 64'b0010100001000000101010101000110110101011010001010000001110010101; end
            14'd3271 : begin out <= 64'b1010101010000111101001000110110010100100000010110001101101000011; end
            14'd3272 : begin out <= 64'b0010100111101001001001110000101100100101000000000010100111101010; end
            14'd3273 : begin out <= 64'b0001110001101010000011011000111010101001111011110001110100111001; end
            14'd3274 : begin out <= 64'b1010100111010001101010011000100000101001110101100010101111010101; end
            14'd3275 : begin out <= 64'b0001011001101101101010011110100100101000001111001010000010000000; end
            14'd3276 : begin out <= 64'b0001110000010001100010111100100010101011010100010010010000000100; end
            14'd3277 : begin out <= 64'b1001101010100010101010001011011110100101010111111010100111000001; end
            14'd3278 : begin out <= 64'b1010011111100000101010001000110110100000110100100010100010010110; end
            14'd3279 : begin out <= 64'b1010101100010000101010000001110000101100001011000001101100100100; end
            14'd3280 : begin out <= 64'b1001101001001100001010101110110100101001101010011010011001101110; end
            14'd3281 : begin out <= 64'b1010000111000111001010001110010010100011110100111010010101000010; end
            14'd3282 : begin out <= 64'b0010000111111010001010110000010100100110110110010010010110101010; end
            14'd3283 : begin out <= 64'b0010100001111010101010000110001000101010000101111010101110001100; end
            14'd3284 : begin out <= 64'b0010000011010011101010010001111110101011011010010001001100010001; end
            14'd3285 : begin out <= 64'b1010100111011111001010101110000000101001100011110010100101001011; end
            14'd3286 : begin out <= 64'b1010010100011110001001110101111110101010111011101010011010111101; end
            14'd3287 : begin out <= 64'b0010100010110111001001101010011010011001101001101010011000101101; end
            14'd3288 : begin out <= 64'b1010010101111010100111101100001100101010101000011010011011010101; end
            14'd3289 : begin out <= 64'b0010010110001111001010001100110100101011110100111010100010101010; end
            14'd3290 : begin out <= 64'b0010101111100100000111101010100100100101011101000010011100001101; end
            14'd3291 : begin out <= 64'b0010100101011000101010001000111110100001111001111010010011101110; end
            14'd3292 : begin out <= 64'b1010101100000100101001101000110110101011011000111010010100010100; end
            14'd3293 : begin out <= 64'b1010100110111100101001001101111010101000010110010010100110010011; end
            14'd3294 : begin out <= 64'b0010000001001111001001110110011110100100010001011010000101111001; end
            14'd3295 : begin out <= 64'b1010100111101111001000000010001000101010101110010010100000111011; end
            14'd3296 : begin out <= 64'b1010101111111110001010000111000110011101110101100010100101000000; end
            14'd3297 : begin out <= 64'b1010100001000011101010000100001010101000000101001010001011010100; end
            14'd3298 : begin out <= 64'b1010100101001011101010111010010010100100110010000010101101100001; end
            14'd3299 : begin out <= 64'b0001000000000111101001001001000010101011001101000001011010110000; end
            14'd3300 : begin out <= 64'b0010100011100001101010111100101010101001100100010001010110110011; end
            14'd3301 : begin out <= 64'b1010101101001011001001100010111100101000000111111010101001000001; end
            14'd3302 : begin out <= 64'b0010100001011011101010101000011000100011010001010010001111101001; end
            14'd3303 : begin out <= 64'b0010011011000110101010011000011000011110000111010010101000011100; end
            14'd3304 : begin out <= 64'b0010101000000111001010000100001010101001110000010010101001011110; end
            14'd3305 : begin out <= 64'b0010101111110111001010101111001100101000111000101010011111110110; end
            14'd3306 : begin out <= 64'b0010011001100001001010111101011000100100101110100010011110101100; end
            14'd3307 : begin out <= 64'b1001110000110000001010100101111010100101101011110001101000011010; end
            14'd3308 : begin out <= 64'b0010100110001100000100100010000110101011000101000010101000110011; end
            14'd3309 : begin out <= 64'b1010011001011011001001001001011100101010011100011010001111001110; end
            14'd3310 : begin out <= 64'b1010100011010011001010001001101000100110011100101010100101110000; end
            14'd3311 : begin out <= 64'b1010010011100100101001111101011110100101100101110010110000101110; end
            14'd3312 : begin out <= 64'b1010011011111001101001000011001010100001110110000001111000100111; end
            14'd3313 : begin out <= 64'b0010010110011000101000111001111010100011000110100010100010010110; end
            14'd3314 : begin out <= 64'b0010100110010010101000010001011110101010000011011001011100111010; end
            14'd3315 : begin out <= 64'b0010101011000100001000101001011110100001101100110010101010101011; end
            14'd3316 : begin out <= 64'b0010100100010100101010111011001100101000011010111001100010011010; end
            14'd3317 : begin out <= 64'b0010101010010110101001011101000100010101000100011010000110000111; end
            14'd3318 : begin out <= 64'b1010011110111011000110111111100010101011001101000001001011011110; end
            14'd3319 : begin out <= 64'b1010100111000111101010100101111100101000000100001010010000110010; end
            14'd3320 : begin out <= 64'b1001101101010111001001110110100110101001110101000010100011111110; end
            14'd3321 : begin out <= 64'b1001111110001001100110011110001000100111010001000010001100000011; end
            14'd3322 : begin out <= 64'b0010010001110111001010000100101100100100101111010010010001110000; end
            14'd3323 : begin out <= 64'b0010011000001011101010101110111000100100111010100010001101001000; end
            14'd3324 : begin out <= 64'b1010100001101000000111101001001110100110001101010010000011000111; end
            14'd3325 : begin out <= 64'b1010011101010000101010010001000100101010011111001010101010000000; end
            14'd3326 : begin out <= 64'b1010100111101111001000001010010110101011001111011010000001110101; end
            14'd3327 : begin out <= 64'b1010001111100101001010101010101100101000011000111010101000010011; end
            14'd3328 : begin out <= 64'b1010011101011010100111010100001010101000110101100010000110100110; end
            14'd3329 : begin out <= 64'b0010100001101011101001011101101010101010111101010010101111101100; end
            14'd3330 : begin out <= 64'b1010101101101000001010100110101110100011100010010010101110111001; end
            14'd3331 : begin out <= 64'b0010101001001010100101110001001100100101010111111010100000001111; end
            14'd3332 : begin out <= 64'b1010100111011101101010110100100000101001100001111010101010001001; end
            14'd3333 : begin out <= 64'b0010101000010110101010101011010010101000100110101010100010100111; end
            14'd3334 : begin out <= 64'b1010100000010001000111110001000100100010100011010010011010011110; end
            14'd3335 : begin out <= 64'b0010010101100111100100011111010110101010010111110010001000100111; end
            14'd3336 : begin out <= 64'b1010000111111111101010101101001110100010110110110010100001110110; end
            14'd3337 : begin out <= 64'b1010010111011100101010110111000100100001000010001010011010010100; end
            14'd3338 : begin out <= 64'b0010010000110111101010010111111000100010100111010010100111000010; end
            14'd3339 : begin out <= 64'b1001110000111001001000001111110010011001011101111010101110100101; end
            14'd3340 : begin out <= 64'b1010100010111110001001111011000110101001010100101010100101111011; end
            14'd3341 : begin out <= 64'b0010100011110011001000001100100010010110000110101010001110100111; end
            14'd3342 : begin out <= 64'b1010001100000111001001011111110010100100011001011010011110101010; end
            14'd3343 : begin out <= 64'b1010010011010111101001110110100100011010111110111010101100010000; end
            14'd3344 : begin out <= 64'b1001100111111111001001110010111100100101000101101010100111110010; end
            14'd3345 : begin out <= 64'b0010101000001100001010100001111000101011000010011010001110011001; end
            14'd3346 : begin out <= 64'b1010011001010000001001010110101110101001000000000010001001011001; end
            14'd3347 : begin out <= 64'b1010100100100000001010100000110100011111001110010010010011110110; end
            14'd3348 : begin out <= 64'b0010010100000001000101000101010100100001011110111010101011100100; end
            14'd3349 : begin out <= 64'b0010001110100001101000011100001100101010011111000010011111100010; end
            14'd3350 : begin out <= 64'b0010000101000101000111010101101010101100000001010010100101010010; end
            14'd3351 : begin out <= 64'b0010001001110111001010110010110110101000110100011001111000111111; end
            14'd3352 : begin out <= 64'b0010101111011010001010001010010110100101110110111010001010000001; end
            14'd3353 : begin out <= 64'b1010101001101111101010001111001000101010101011100010101011101010; end
            14'd3354 : begin out <= 64'b1010100100011001101001101001100010100110000010000001100000010110; end
            14'd3355 : begin out <= 64'b0010010011110100001010101011010110101011010010000001101110000000; end
            14'd3356 : begin out <= 64'b0010100100010111101010011101100010101000110011100010100001010000; end
            14'd3357 : begin out <= 64'b1001111111011001001000100011100010001010100110000010010010111001; end
            14'd3358 : begin out <= 64'b1001110011100100100111011101000010100010010101001010100000010100; end
            14'd3359 : begin out <= 64'b0010101101001010101010111100000100100100010110110010011110100010; end
            14'd3360 : begin out <= 64'b1010011111110000001010011111011010101011000001111010010001010110; end
            14'd3361 : begin out <= 64'b1010100110011111101010111111111110101010000100010010010111001110; end
            14'd3362 : begin out <= 64'b0010001000100010001001011110111010100011001110010010100010101101; end
            14'd3363 : begin out <= 64'b0010101111010010101010010111000010101010001001001010101011010110; end
            14'd3364 : begin out <= 64'b0010010111011110001001011111101110100001011010010010100000101111; end
            14'd3365 : begin out <= 64'b1010101111001000100111100000001110100101010110101010101001010110; end
            14'd3366 : begin out <= 64'b1001111011110110000101100011110000101000101000100010100000111010; end
            14'd3367 : begin out <= 64'b1010101000011111001000100010111100101001001001111001110001100110; end
            14'd3368 : begin out <= 64'b1010101110010111001001010011111010101011001111001010100100101010; end
            14'd3369 : begin out <= 64'b1010000110000010101010101011101010011101101110100010100110010100; end
            14'd3370 : begin out <= 64'b1010011000010111000011010111001110101000110100001001100110110000; end
            14'd3371 : begin out <= 64'b1010101000110110001010111100000100011011011011100010011100101101; end
            14'd3372 : begin out <= 64'b0010110000010111001010100101001100101001111010111010010101101010; end
            14'd3373 : begin out <= 64'b1010000101001001101010000100100000101000000001010010100010101101; end
            14'd3374 : begin out <= 64'b0010000100000010100111110001011100101000000000011010100010001010; end
            14'd3375 : begin out <= 64'b0010100010110111101000000100111000101001011111101010011000000001; end
            14'd3376 : begin out <= 64'b1010010011010010001000010111111110100100111000001010010000000011; end
            14'd3377 : begin out <= 64'b0010011001011011101001011101000000100111000000111001001001010111; end
            14'd3378 : begin out <= 64'b1001110111110000001001000000010100101000101000000010010001101100; end
            14'd3379 : begin out <= 64'b1010100000110001101010100110011100100110110001110010100110010011; end
            14'd3380 : begin out <= 64'b1010100111010001101010001000101000100100101001111010011100000100; end
            14'd3381 : begin out <= 64'b1010101100001011001010001000110100101010100000111010011000111001; end
            14'd3382 : begin out <= 64'b0010010110011001101000111101101100101011110101110010100110011000; end
            14'd3383 : begin out <= 64'b1010001111010011001010001010001000100101110100110010010100011100; end
            14'd3384 : begin out <= 64'b0010001101001000000111010000010110100111001110000010000100000000; end
            14'd3385 : begin out <= 64'b0010000101100000100110100010010010100100000001110010000010110110; end
            14'd3386 : begin out <= 64'b1010101100001110101001010110001100101010011000000010000010110001; end
            14'd3387 : begin out <= 64'b1010100010101110001000101101110000101011101101100010100111110011; end
            14'd3388 : begin out <= 64'b0010101011010000001000110011010010101011111001010010101001111001; end
            14'd3389 : begin out <= 64'b1010011100011111101000011111111100101001100011111010010110000001; end
            14'd3390 : begin out <= 64'b1010010101101100001001100101110100100110001000010010101000011010; end
            14'd3391 : begin out <= 64'b1010100011111100101000000010010110101001101111111010101001011010; end
            14'd3392 : begin out <= 64'b0010101110010101001000001001011000011111011110011010101010001101; end
            14'd3393 : begin out <= 64'b1010001000100100101010110010011010101001010111101010000000001000; end
            14'd3394 : begin out <= 64'b0010000110000000001010100001110110101010100011111010100100010000; end
            14'd3395 : begin out <= 64'b1010110000100101100111010100010100011101010111111010100101111001; end
            14'd3396 : begin out <= 64'b1010101100101011101000101001000100101010101011101010001001000001; end
            14'd3397 : begin out <= 64'b1010101100101000001010011001101110100100011010011010000100100110; end
            14'd3398 : begin out <= 64'b0010101001111010001010011000101000100111000110011010001001000111; end
            14'd3399 : begin out <= 64'b0010101101001101000111100010100110101011011010000010001101010100; end
            14'd3400 : begin out <= 64'b1010100100000011101000000111110110010111100111010010010001000110; end
            14'd3401 : begin out <= 64'b1010011110110000001001000000010010010101001110010010101001011110; end
            14'd3402 : begin out <= 64'b0010100011011100001001001101001010100010000110011010110001000101; end
            14'd3403 : begin out <= 64'b0010101010100100001001110100111100101000100100110010101110010101; end
            14'd3404 : begin out <= 64'b1001100011011001100111001011011100100100000011010010101101111100; end
            14'd3405 : begin out <= 64'b1000111101000100101010110101011100100110101111001010101100100101; end
            14'd3406 : begin out <= 64'b1010011000101101101000010001110000100111010000010010000111010000; end
            14'd3407 : begin out <= 64'b0010010000101111101010010011010100101010011000111001100100100101; end
            14'd3408 : begin out <= 64'b1010101000000000101010011010100010100011100100100010101110001011; end
            14'd3409 : begin out <= 64'b0010101100111000001010110001000010100101100010101010010010001000; end
            14'd3410 : begin out <= 64'b0010101011010001000110000111011010100010000101111010101110110010; end
            14'd3411 : begin out <= 64'b1010101101011101001010111100001100100000111010101010100010111011; end
            14'd3412 : begin out <= 64'b0010010101011111101000100000100010101001000010111010100011000111; end
            14'd3413 : begin out <= 64'b0010100100110100101010010001000100100010011010010001101110010110; end
            14'd3414 : begin out <= 64'b0010101001010110101001111011011100100000000000111010101110011010; end
            14'd3415 : begin out <= 64'b1010100011001001101010000110010100100100101001010010000000001100; end
            14'd3416 : begin out <= 64'b1010010000100011101001101111111000100110001011010010101111010101; end
            14'd3417 : begin out <= 64'b1010000110101100100110001111001010101100000101100010100100010000; end
            14'd3418 : begin out <= 64'b1001111011110110001001010101001110101001111010110010100110000101; end
            14'd3419 : begin out <= 64'b1010100110100101001000001000110100101000111111001010101100011101; end
            14'd3420 : begin out <= 64'b0001101000010111001001101101101000100100100111100010101011011011; end
            14'd3421 : begin out <= 64'b1010011110011010101001101001000110100001010111111010101000000001; end
            14'd3422 : begin out <= 64'b1010101100010101001010011111000010011010000110100010101011111010; end
            14'd3423 : begin out <= 64'b0001101011000011101010001111101000100000010100110010001110101000; end
            14'd3424 : begin out <= 64'b0010101010100101101001001111011000101001010011010010011100111101; end
            14'd3425 : begin out <= 64'b0010100000011001101010011001101010101000011000111001111100100100; end
            14'd3426 : begin out <= 64'b0010011011001001001001001000010110100011011101100010101111000011; end
            14'd3427 : begin out <= 64'b0010100111000111000100110000011010100101100011111010100100011011; end
            14'd3428 : begin out <= 64'b1001100100101101101010010110001110011100000011001010100011110001; end
            14'd3429 : begin out <= 64'b0010101100111100001010011010111010101001010010100010101100111011; end
            14'd3430 : begin out <= 64'b0010101001011110001001111000011100101010111100010001101001110110; end
            14'd3431 : begin out <= 64'b1010010000001101101001110001001110100100111100011010010110011101; end
            14'd3432 : begin out <= 64'b0001110110100011101010110101111000101000011101100010100100011011; end
            14'd3433 : begin out <= 64'b1010101000001011001010000101100010101001100001101010101001010100; end
            14'd3434 : begin out <= 64'b0010011110100010101010010000010000100000110111101010001000100001; end
            14'd3435 : begin out <= 64'b0010011000100110001010000111100110100011011001000010101101010011; end
            14'd3436 : begin out <= 64'b1010101111111111101010110110011100100101111010000010010010101010; end
            14'd3437 : begin out <= 64'b0001101011100010000111000011000110101000111100000010001100101001; end
            14'd3438 : begin out <= 64'b1010101001100111001010110100011100101010100110010010101000011100; end
            14'd3439 : begin out <= 64'b0010000101011101000111110101111110100111111001110010101000101011; end
            14'd3440 : begin out <= 64'b0010100111010011001010101111000110101001010011010010011000110100; end
            14'd3441 : begin out <= 64'b0010011011001101101010010101001110101010011110010010010111110100; end
            14'd3442 : begin out <= 64'b1010100111100011001010010010000100100110110001011010101011101010; end
            14'd3443 : begin out <= 64'b1010101011011100001001100010000000101000111010111001101011111001; end
            14'd3444 : begin out <= 64'b0010100111101101101001001111100110010101000101010010100100100011; end
            14'd3445 : begin out <= 64'b1010010010100101101000010011110110101000011001001001111110110001; end
            14'd3446 : begin out <= 64'b0001111001101010001001010010001110101010110101011001011001110110; end
            14'd3447 : begin out <= 64'b0010110001010011101010001000110000100110101101110010100001001100; end
            14'd3448 : begin out <= 64'b1010000000011111001010010111000110101001011001010010000100100000; end
            14'd3449 : begin out <= 64'b1001001111010101000111101101011110100110111111010010100101010000; end
            14'd3450 : begin out <= 64'b0010001110111000101010111111111110101000010010001010101100101010; end
            14'd3451 : begin out <= 64'b0010100000011100001000100100100110100011010001011010001101100010; end
            14'd3452 : begin out <= 64'b0010100000000110101010001101111010101011110000000010010010100111; end
            14'd3453 : begin out <= 64'b1001111010101110101010110111000000101000010110001001111100000101; end
            14'd3454 : begin out <= 64'b0010101110101011101010110111111100100110001110101010100011101000; end
            14'd3455 : begin out <= 64'b0010000110011111101010001110110000101010111101100010100010000010; end
            14'd3456 : begin out <= 64'b0010101110010001001000011111111010100100010101101010101111111011; end
            14'd3457 : begin out <= 64'b0010101000000011001001011001100010101000100100011001100011101010; end
            14'd3458 : begin out <= 64'b1010100010011110001001111110011100101010101110001010010010010001; end
            14'd3459 : begin out <= 64'b1000110111100001001010001011111000101000001110001010101001101001; end
            14'd3460 : begin out <= 64'b0010100100101100101010110001100000100000001010011010100011010111; end
            14'd3461 : begin out <= 64'b0010000111011010001001110111011010101001011000000010110000010001; end
            14'd3462 : begin out <= 64'b0010011001010000001001111001011000101000101110011001011100101001; end
            14'd3463 : begin out <= 64'b0010011100000101101010000110010110100000100111100010010000010010; end
            14'd3464 : begin out <= 64'b0010101110000010001010111100011100101010000011000010010000110010; end
            14'd3465 : begin out <= 64'b1010000111001000001000011110101100101001001100101010001110000110; end
            14'd3466 : begin out <= 64'b0001011111010001001010110110011110101011101011110000101101010001; end
            14'd3467 : begin out <= 64'b0010100100011110001010011110100110101001011110001010010101110111; end
            14'd3468 : begin out <= 64'b1010101011101101100100111010101000101011111100100010100110011001; end
            14'd3469 : begin out <= 64'b1010001000011001101000100101111100101010011011111010101111000100; end
            14'd3470 : begin out <= 64'b0010010110001100101010111010101010100110010000000010101011001010; end
            14'd3471 : begin out <= 64'b1010011011001010001010100001100100101011011001001010101010001010; end
            14'd3472 : begin out <= 64'b0010011011101110001001110011110000101001000001010010100000000101; end
            14'd3473 : begin out <= 64'b0010100111001111101001011011000000101010001111111010010000110001; end
            14'd3474 : begin out <= 64'b1010011110010010001001100101011010100111011101010010000111001001; end
            14'd3475 : begin out <= 64'b0010100110110000100110110100011010101011010011001001101111111000; end
            14'd3476 : begin out <= 64'b0010100111101001001000111110101100101001010110110010101111011000; end
            14'd3477 : begin out <= 64'b1000111100100111001000011100011100101000001110110010101110010111; end
            14'd3478 : begin out <= 64'b0010001010101011001010011100111110101001101011101010100100101011; end
            14'd3479 : begin out <= 64'b0010100001100100101010000001010110100111100100001001100001001001; end
            14'd3480 : begin out <= 64'b0001011001111100001010000101111010101011101010010001011010101001; end
            14'd3481 : begin out <= 64'b0010101101011111000111001001000110101001111100100001111101000101; end
            14'd3482 : begin out <= 64'b0010101001101111001000000001000100101000101111101001111011111001; end
            14'd3483 : begin out <= 64'b1010100111000110001010110010101000100111001000010010010010110001; end
            14'd3484 : begin out <= 64'b1010101001111100101001110000101010101010011011000010010010111011; end
            14'd3485 : begin out <= 64'b0010010001100101100111000111100010101001110111110010101111010101; end
            14'd3486 : begin out <= 64'b1010100100100000001010101101010100101000010010000010011110011010; end
            14'd3487 : begin out <= 64'b1010011100110110101010111100011000100111100011011010101101111000; end
            14'd3488 : begin out <= 64'b1010101000001011001010100101001000100001011100001010100100010100; end
            14'd3489 : begin out <= 64'b0010000010110011101010010101111010100010110000101001111010000100; end
            14'd3490 : begin out <= 64'b1010100010100100101010011101010000100111101101100001111010101000; end
            14'd3491 : begin out <= 64'b1010000001100010101001000001010010101000110001010010101010011100; end
            14'd3492 : begin out <= 64'b0010100010110011001010001011001010100000111111000010011000101100; end
            14'd3493 : begin out <= 64'b0010100111001110001000010010000010100011111111011010011011000100; end
            14'd3494 : begin out <= 64'b1010000001010111001010100011001000100101001001011010100011010100; end
            14'd3495 : begin out <= 64'b0010101000111000101001000001000110101010001010111010010001110110; end
            14'd3496 : begin out <= 64'b1010010101011111001010110111101110101000000010010010100010110000; end
            14'd3497 : begin out <= 64'b1010000010001001001001010010000000101010011111000010101100011111; end
            14'd3498 : begin out <= 64'b0010101000100011001000011101010010101011111111011010101111000011; end
            14'd3499 : begin out <= 64'b0010101000111001101010100100000100010110010001111001010010110111; end
            14'd3500 : begin out <= 64'b0010010000011111101010111101101000100110001110001010100110111100; end
            14'd3501 : begin out <= 64'b0010100110110100001001100111011110100111101101110001100010011100; end
            14'd3502 : begin out <= 64'b0010101111011010101010010011010000101001000101110010100000101010; end
            14'd3503 : begin out <= 64'b0010010001100011000110101010011010100100110100001010100001011001; end
            14'd3504 : begin out <= 64'b1010000001010100101001110101011010101011010100101010100001010100; end
            14'd3505 : begin out <= 64'b1010011100001000101001010000100010010101101110111010100011010001; end
            14'd3506 : begin out <= 64'b0010100111010011100111101001111110101001001110100010110000011011; end
            14'd3507 : begin out <= 64'b0010100001110000101001101100011110101001001011100010100010100001; end
            14'd3508 : begin out <= 64'b1010101011101011101010111000111000011110011010001001101110101010; end
            14'd3509 : begin out <= 64'b1010101110000111101001111100101110100111001001101001111101011101; end
            14'd3510 : begin out <= 64'b0010101010011011001000000011011000100011111100101010010010100010; end
            14'd3511 : begin out <= 64'b1010011001001001101001011000001000101000011100110010101010000101; end
            14'd3512 : begin out <= 64'b0010011000000110100101111010010000100101010110111010101001100010; end
            14'd3513 : begin out <= 64'b0010011010101001001001001110011000101010011111010010011000101010; end
            14'd3514 : begin out <= 64'b0010011011100101001001111111001100100111000000110010011100101000; end
            14'd3515 : begin out <= 64'b0010110001001000101010101110010010100100010001100010010011110110; end
            14'd3516 : begin out <= 64'b0010100000011111000101000101011110100010101000001010010101110101; end
            14'd3517 : begin out <= 64'b1010000000011010001010011101010100100110011100111010110000001110; end
            14'd3518 : begin out <= 64'b0010101100100000101000100100000000100101011010101010100000111101; end
            14'd3519 : begin out <= 64'b1010000100101101101010100001000110101010100011111010100010100110; end
            14'd3520 : begin out <= 64'b0010101011100100000111100000011110101011110000001010100011110100; end
            14'd3521 : begin out <= 64'b0010100110011100001010110100101000101010001000101001110111000011; end
            14'd3522 : begin out <= 64'b1010000101110100101001101010110100100101001101110010000101010011; end
            14'd3523 : begin out <= 64'b1010101110101100001001110100110100100011000001110010101010000000; end
            14'd3524 : begin out <= 64'b0001111011101111001001101010011000100110100010000010010010100000; end
            14'd3525 : begin out <= 64'b1010101000001001101010010011111000101011000101101001110101101111; end
            14'd3526 : begin out <= 64'b1010011110111100101010010011101100100101100111011010010100000110; end
            14'd3527 : begin out <= 64'b1010101100111001001000001011011110101011001101010010101110011000; end
            14'd3528 : begin out <= 64'b0010100001101101001010111111011100100100000101000010101101000000; end
            14'd3529 : begin out <= 64'b1010100101110101101010011100010000011111011111010010101110010001; end
            14'd3530 : begin out <= 64'b0010010001110100001010111111001010100011110011111010100010011010; end
            14'd3531 : begin out <= 64'b0010101111000110001001101101111110101001010110100010100100000100; end
            14'd3532 : begin out <= 64'b1010010100000110001001011101010010100010111011101010001001111011; end
            14'd3533 : begin out <= 64'b0010011111110011101010001011000010101010111001100010001101000101; end
            14'd3534 : begin out <= 64'b1010000101101011101001001111011000101011101001111010101110011011; end
            14'd3535 : begin out <= 64'b1001101001000111101010111001001000101011010100110010101111001000; end
            14'd3536 : begin out <= 64'b0010100001100010001010111001101000101000001000010010010101100011; end
            14'd3537 : begin out <= 64'b1010000011000101000100111011000110100111010011101010100011111110; end
            14'd3538 : begin out <= 64'b0010101100110110001010011111100010101000000101000010110001000001; end
            14'd3539 : begin out <= 64'b1010010011111110101010001101101110101010100100001010101111100010; end
            14'd3540 : begin out <= 64'b1010101011111001000111110001110100101010101110000010011000100010; end
            14'd3541 : begin out <= 64'b0010001011101110101000001110111110100111011111000001011010010000; end
            14'd3542 : begin out <= 64'b0010011110010011001000111000000000100111011111110010001000010111; end
            14'd3543 : begin out <= 64'b0000101110110011101010100000000010101001111100101010001101111111; end
            14'd3544 : begin out <= 64'b1010000000010111001001110011011010101001110011000010101100101110; end
            14'd3545 : begin out <= 64'b0010101011110011101010001011000010100100100001100010100011001111; end
            14'd3546 : begin out <= 64'b1010100110001101101010000000110010101010001111010001010101110000; end
            14'd3547 : begin out <= 64'b1010100100110101101001111010111110101001111111001010010110010100; end
            14'd3548 : begin out <= 64'b0010010011000010101001100110011110101000101011100010100110011101; end
            14'd3549 : begin out <= 64'b1001101111100110001010010100100010101000001100111010101010111101; end
            14'd3550 : begin out <= 64'b1010101011110011001010011110001010011111101100111010000110111000; end
            14'd3551 : begin out <= 64'b0010010100001011101010100000100000000001110011110001111001100011; end
            14'd3552 : begin out <= 64'b0010000000100111101010011110010100011100000100100010100100000011; end
            14'd3553 : begin out <= 64'b0010000001111001101001010011110000101001010110000010010011000000; end
            14'd3554 : begin out <= 64'b1010100011111001101010001010100110100100011110010010101101011100; end
            14'd3555 : begin out <= 64'b1010000000011110101010000010100110100001010010111010100001110011; end
            14'd3556 : begin out <= 64'b0010000011000001001001010011001000101001001100000001011011010000; end
            14'd3557 : begin out <= 64'b0010100101100001001001010111011000101010010101111001111110001001; end
            14'd3558 : begin out <= 64'b1010101000010011100110100011000110100110001001101010010101000000; end
            14'd3559 : begin out <= 64'b0010011010000001101001100010001100000011001110100001110010101010; end
            14'd3560 : begin out <= 64'b0010000111100111001010100001101110101010000110011010100001001011; end
            14'd3561 : begin out <= 64'b1010011001110110001001110000001000101001000101000010101110101001; end
            14'd3562 : begin out <= 64'b0010100100010100101010001101111010100101111001101010100001111100; end
            14'd3563 : begin out <= 64'b0010001010101110101000100010111000100010101001100010100101100100; end
            14'd3564 : begin out <= 64'b1000011110011001001010110110011110101000100001001010001000100101; end
            14'd3565 : begin out <= 64'b0010101011111001101000000110011000011110101001100010010010011110; end
            14'd3566 : begin out <= 64'b1010100001111011001010011101011010101001101101111001110001101111; end
            14'd3567 : begin out <= 64'b0010101011110100000111001110111110101011100100111010101100101000; end
            14'd3568 : begin out <= 64'b1010101100010001101010110101011010101011111101101010101111101101; end
            14'd3569 : begin out <= 64'b0001010101000100000110100001001000101001111000101010101110101110; end
            14'd3570 : begin out <= 64'b1010011101000110101010111101100010101011101110111010010001110010; end
            14'd3571 : begin out <= 64'b0010101010100001101010100000000010101011011011110010010100011001; end
            14'd3572 : begin out <= 64'b0010000100011001101010000100000010100110011101010010001011110100; end
            14'd3573 : begin out <= 64'b1010101011001100001001110001100110101010101000011010011100001100; end
            14'd3574 : begin out <= 64'b1010101101001101101010001001101000101000011011110010100001101010; end
            14'd3575 : begin out <= 64'b1010101000010111001010011110100100101000100100111010000100010000; end
            14'd3576 : begin out <= 64'b1010010010011011001001101011110000101010001100001010011100100010; end
            14'd3577 : begin out <= 64'b0010011100110010001010111001011000100010111100010010010100111100; end
            14'd3578 : begin out <= 64'b1001011101111110101000101011100100101001111010110010000000101101; end
            14'd3579 : begin out <= 64'b1010101010010001101010111010110010101011010100110010101000010110; end
            14'd3580 : begin out <= 64'b1001101110111011101010111011000110100101111011010010000110101000; end
            14'd3581 : begin out <= 64'b0010001011101110001010001001000100101011100100010001010100110100; end
            14'd3582 : begin out <= 64'b1010100110000000100110111101010100101000011100011001011100110011; end
            14'd3583 : begin out <= 64'b0010001010001110101001110011011010100000100011011010100101011110; end
            14'd3584 : begin out <= 64'b0010001001011000100111000011000100101010011110011001111001011100; end
            14'd3585 : begin out <= 64'b0010001001110000001000110100010110101010111000111001101001001000; end
            14'd3586 : begin out <= 64'b1001111111111101101001101010000000101011010010100010101001110001; end
            14'd3587 : begin out <= 64'b0001010000000010001000011110110110100110111001000010011011010101; end
            14'd3588 : begin out <= 64'b0010010001101011101010100110111100100111010011001010011011010101; end
            14'd3589 : begin out <= 64'b0010000100100101101001100001000110100100001010110010100011011011; end
            14'd3590 : begin out <= 64'b0010101111101001001010001101000010100001110110010010100011000001; end
            14'd3591 : begin out <= 64'b1001110010010110101001001011101110101010001101110010010000010100; end
            14'd3592 : begin out <= 64'b1010100111110011100100011000001010011111101100010010001010110010; end
            14'd3593 : begin out <= 64'b0010101100010001001001001011110010101010010100001010101001100110; end
            14'd3594 : begin out <= 64'b0010010000001101101000111001110110100101111111110010101000010110; end
            14'd3595 : begin out <= 64'b1001010000000101101010000110101100101011011000100010010011111000; end
            14'd3596 : begin out <= 64'b1010011001111001001010101011000100100100011011100010100111101101; end
            14'd3597 : begin out <= 64'b0010001100000010000110101010010010101001011111000010101011111110; end
            14'd3598 : begin out <= 64'b1001111000000011101000100011110010100101111000111010101101000000; end
            14'd3599 : begin out <= 64'b1010100111111010001010011110001100100001000101100010100111100000; end
            14'd3600 : begin out <= 64'b1010001110010111101010011100011110101011101010111001111100111101; end
            14'd3601 : begin out <= 64'b0010000001100011001000011111110100011010010111010010100110000011; end
            14'd3602 : begin out <= 64'b1001100101001000001010001010101010100001111011010010001010110100; end
            14'd3603 : begin out <= 64'b1010101001100000001001011100111000010101110111001010000100111000; end
            14'd3604 : begin out <= 64'b0010010000000111001001010000111110100100011000010010000001010011; end
            14'd3605 : begin out <= 64'b1010100001111100101010001100001110100010100111111010011101010101; end
            14'd3606 : begin out <= 64'b1000111000000100001010000111101010101100000010000010101011101111; end
            14'd3607 : begin out <= 64'b1010101000100110101010111010111000101001000011101010101110011100; end
            14'd3608 : begin out <= 64'b1010101000001101101010001100110010101001110000101001100011000000; end
            14'd3609 : begin out <= 64'b0010100110101001001010001100001100101001100101011010100001110111; end
            14'd3610 : begin out <= 64'b0010011101110011101010101101111000101001101000010010100100100100; end
            14'd3611 : begin out <= 64'b0010101001001110101010001100100000100100011001001010001111111101; end
            14'd3612 : begin out <= 64'b1010100100110001000111001100111110101011000010100010010011100010; end
            14'd3613 : begin out <= 64'b0000011100110110001010110110100000101000110111110010000011000101; end
            14'd3614 : begin out <= 64'b0010101100010001101010100101101110101011000110110010000010110100; end
            14'd3615 : begin out <= 64'b0010010010110011101001100010100100101011100111111010101100010111; end
            14'd3616 : begin out <= 64'b0010011010011101101001010000001000100010111101011010100110101111; end
            14'd3617 : begin out <= 64'b1010100000101100101000111011110000011110001000101010010001011100; end
            14'd3618 : begin out <= 64'b0010101001001010101010000011000100101000011111010010100111010100; end
            14'd3619 : begin out <= 64'b0010001110101001001000001111001010100101110111001010100000011011; end
            14'd3620 : begin out <= 64'b1010110000001100101010110010011110101010101101110010010010111001; end
            14'd3621 : begin out <= 64'b0010011101011010001010011001100100101010100011110010101011011010; end
            14'd3622 : begin out <= 64'b1010001100110010001010000010010000101001011001111010011001011110; end
            14'd3623 : begin out <= 64'b1010011100110001001000000011010000011110000001110010101000111100; end
            14'd3624 : begin out <= 64'b0010011100011111001010010110010110101000010111010010100111100100; end
            14'd3625 : begin out <= 64'b1001100101001110101010000110011110101001110000101010100000101110; end
            14'd3626 : begin out <= 64'b1010100101111001101010010000011000100011011011101010101111100100; end
            14'd3627 : begin out <= 64'b1010001010111110101001001110110010101011001000010010100100100001; end
            14'd3628 : begin out <= 64'b0010100000111011101001111000010100011010110011000010100101110100; end
            14'd3629 : begin out <= 64'b0010100001001000101000100010101000100110001111001010011010100001; end
            14'd3630 : begin out <= 64'b0010100100110100001010010010000100101001011111010010000010101011; end
            14'd3631 : begin out <= 64'b1010000011000001001001110000111000100101100110110010011011111001; end
            14'd3632 : begin out <= 64'b1010011110111011100101110010110010100110100001101010101000001010; end
            14'd3633 : begin out <= 64'b1010101011110010101001000001101010010111110100000010100100000101; end
            14'd3634 : begin out <= 64'b0001100100000100001000111001001000101001101000010010100001001101; end
            14'd3635 : begin out <= 64'b0010100101100101001001100001100010101011111101001010010101010000; end
            14'd3636 : begin out <= 64'b0010100001110110101000011101100010011110001001010010000000110110; end
            14'd3637 : begin out <= 64'b1010101010101011001010110111100100101001110011000010101011011100; end
            14'd3638 : begin out <= 64'b1001110101100010101010111110111110101001110010100010011001010110; end
            14'd3639 : begin out <= 64'b1010100110010001000101000000011010101000110010101010010001001110; end
            14'd3640 : begin out <= 64'b1010010110101011001010101101101110101010100110010010001001111001; end
            14'd3641 : begin out <= 64'b1010011000011100101000001010010010100011101011000010100011001100; end
            14'd3642 : begin out <= 64'b1010000000001101101000000001001100100001010111111010101000011010; end
            14'd3643 : begin out <= 64'b0010101011100111101001110100010110100111010011000001100011101000; end
            14'd3644 : begin out <= 64'b0001101010110111001001101011101000010100010100110010101110000000; end
            14'd3645 : begin out <= 64'b1010011100101101100111100111000000101011010001000010101110111110; end
            14'd3646 : begin out <= 64'b0001110100100100101000010110110000101000011000011010101001000010; end
            14'd3647 : begin out <= 64'b0010011111010010101010000000011000100101000010001010100001010111; end
            14'd3648 : begin out <= 64'b0010100110001011101010101011010110101010001000101010011010111111; end
            14'd3649 : begin out <= 64'b0001111110011011101010010101110100011100011110000010100011110101; end
            14'd3650 : begin out <= 64'b1010100011000011101000011010010010101011000000001010101100110111; end
            14'd3651 : begin out <= 64'b1010101100110011100110111010000010100101111100111010100111100010; end
            14'd3652 : begin out <= 64'b0010001001111100101010100110000100101011111110110001110011100001; end
            14'd3653 : begin out <= 64'b0010101110000110100111100001100110101010011011111010100101110000; end
            14'd3654 : begin out <= 64'b1001110010100010001000111011101100101010011110000010100011001010; end
            14'd3655 : begin out <= 64'b0010010100000111001001100110001100100101110000110010100100100111; end
            14'd3656 : begin out <= 64'b0001111100010110001010101011010010101011000001110010101110000011; end
            14'd3657 : begin out <= 64'b1010001011000111001010001100110100101010101110100010100111100011; end
            14'd3658 : begin out <= 64'b0010000111000011001010110100110000100100110100100010001101110000; end
            14'd3659 : begin out <= 64'b0010101010111111101000101100110100100111010101010010011000000010; end
            14'd3660 : begin out <= 64'b0001100111001011001001111100010010101010100010111010011100010000; end
            14'd3661 : begin out <= 64'b0010101111000111101010101011110110010001101000100001000111001010; end
            14'd3662 : begin out <= 64'b1010100100100011101010100001100010101011011110001010001110000010; end
            14'd3663 : begin out <= 64'b1001110101000000101010101110001010100101100011111010101101000001; end
            14'd3664 : begin out <= 64'b0010010101111110001000000101100010101011111000000010100110000000; end
            14'd3665 : begin out <= 64'b1010010000010110101001001100110010101001101011010010011010101110; end
            14'd3666 : begin out <= 64'b0010011011101100101010111011010010100000001010011010011000100001; end
            14'd3667 : begin out <= 64'b1000001110110001100110010110101110101001011011010010100011010011; end
            14'd3668 : begin out <= 64'b1001110000010010101010001010010000100011111000111010000101010010; end
            14'd3669 : begin out <= 64'b1010000010101101100110110010000000100101101111101010010011011100; end
            14'd3670 : begin out <= 64'b1010101100110111101010011000110110101000011010011010001011000001; end
            14'd3671 : begin out <= 64'b0001000111100011001010101111001110100100011010010010010001011101; end
            14'd3672 : begin out <= 64'b0010101000011010001000100001010010101001101110000010010011100110; end
            14'd3673 : begin out <= 64'b0010101000000101001010001010011110100101010111110001011101110010; end
            14'd3674 : begin out <= 64'b0010101010100010101010101001001100101001100011111001110110010000; end
            14'd3675 : begin out <= 64'b0010100010011110100100001110101010101000101001001010010110101011; end
            14'd3676 : begin out <= 64'b1010011001101010001011000100101100101011110111100010100010000010; end
            14'd3677 : begin out <= 64'b1010011001100000101010111100101010100000101011111010011001101100; end
            14'd3678 : begin out <= 64'b0010000110110010001001110001110110101001110001100010101111011110; end
            14'd3679 : begin out <= 64'b0010010100101111100111101110000010100000011101001010101111001010; end
            14'd3680 : begin out <= 64'b1010101110000111101001100010010100100111000100110010100010100010; end
            14'd3681 : begin out <= 64'b1010011111111001001000100110001100101010011010100010010000110001; end
            14'd3682 : begin out <= 64'b1001111100000100101001111101000100101001010001011010100111100110; end
            14'd3683 : begin out <= 64'b1010010011000100101010110111101100101010010010011010100010001100; end
            14'd3684 : begin out <= 64'b0001010110001010101000111110011100101000000110010010100100010010; end
            14'd3685 : begin out <= 64'b1001101110000110001010011000001110011110010110100010101010010101; end
            14'd3686 : begin out <= 64'b1010101101000111000100101110110100100100110110100010011100010101; end
            14'd3687 : begin out <= 64'b1010010111110000101001010011110000011110101111010010101101011010; end
            14'd3688 : begin out <= 64'b0010100110000010001001001101010100101011000011011010100100000000; end
            14'd3689 : begin out <= 64'b1001110111110110101001101100110010101010001111100010010001001000; end
            14'd3690 : begin out <= 64'b0010011101001011001010000101111110101000111100100010011000010100; end
            14'd3691 : begin out <= 64'b0010100011101011001010100101001010101010001000000010000110011101; end
            14'd3692 : begin out <= 64'b0010010111110001000111111011011110100101000110010010011010001101; end
            14'd3693 : begin out <= 64'b0010011101100110101010110011001100100111001110011010100100011100; end
            14'd3694 : begin out <= 64'b0010011101111010100101011010100100101010100001001001111100110111; end
            14'd3695 : begin out <= 64'b1010100001001000100100111100011110100111011100001010011100010110; end
            14'd3696 : begin out <= 64'b0010100111000010001011000010101010101011111000100010101001000110; end
            14'd3697 : begin out <= 64'b1001111000010100001010010011111110100111011001011010101111011101; end
            14'd3698 : begin out <= 64'b1010010001100101101001101100001000100010000101101010000110111010; end
            14'd3699 : begin out <= 64'b0010100011101111001010001100010110010100001101100010011110110100; end
            14'd3700 : begin out <= 64'b0010100100010001000110001001010010011100100001001010000100100001; end
            14'd3701 : begin out <= 64'b0010101111110000101001111010111010100110011010111010010110011011; end
            14'd3702 : begin out <= 64'b1010101000111111101010011011001110100110100100111010101001110110; end
            14'd3703 : begin out <= 64'b0001111010010010001001101001110110101000100101100010010010110110; end
            14'd3704 : begin out <= 64'b0010100101111000101001111000100000101000111000101010101111100001; end
            14'd3705 : begin out <= 64'b0010011100010001101010101011010100100011000001010010000100100110; end
            14'd3706 : begin out <= 64'b1010101011100111001010011010110000101011001110010010011011100110; end
            14'd3707 : begin out <= 64'b0010100100011011001000110001001000101000101101111010100000010101; end
            14'd3708 : begin out <= 64'b0001001110010000001000110001010100101011101011000010010100001011; end
            14'd3709 : begin out <= 64'b0010100100100101101010010001110010100111100110110010100100010011; end
            14'd3710 : begin out <= 64'b0001110101001001100111011110011010101000110000110010100110010111; end
            14'd3711 : begin out <= 64'b1010100111000101001011000001000100001101110001110010100101101010; end
            14'd3712 : begin out <= 64'b1001101001110000101010001000000010100010010011011010100111110110; end
            14'd3713 : begin out <= 64'b0010010101110000101000111110100100011011110110101001110010000011; end
            14'd3714 : begin out <= 64'b1010101100011101101010111000111000100101111111010010101001011101; end
            14'd3715 : begin out <= 64'b0010010010010010101010000000001110101000011111001010010101110101; end
            14'd3716 : begin out <= 64'b1010101001000101101000111101000000101001001110000001110000000011; end
            14'd3717 : begin out <= 64'b0010101100000000001010101111000110101010110011111010011001101011; end
            14'd3718 : begin out <= 64'b0010011110011100101001101000010010100001011000010010100011001111; end
            14'd3719 : begin out <= 64'b0010011011111000101010010010110000010100100101111010100010100100; end
            14'd3720 : begin out <= 64'b0010011111010001001010101100010110100101100101101010001010010101; end
            14'd3721 : begin out <= 64'b0010100000111111101010000101100110011010010011111010100000000101; end
            14'd3722 : begin out <= 64'b0010101010110000001010111111011000100101000011101010001011010100; end
            14'd3723 : begin out <= 64'b1010100011100101101010000001010100101010100110111010100001001010; end
            14'd3724 : begin out <= 64'b0010101001111100001010110110010110101001110011001010101101000000; end
            14'd3725 : begin out <= 64'b0010010011011110101010100101101010011000110101111010010000111010; end
            14'd3726 : begin out <= 64'b0010011111101100101010101001101110101011100101101001100101000001; end
            14'd3727 : begin out <= 64'b1010100001000000101001100111100010100010010111100010001011101111; end
            14'd3728 : begin out <= 64'b0000101010001101101000011011100100101010100110010010100111011100; end
            14'd3729 : begin out <= 64'b1010101001000100101000001010111000010110101111001010101110100001; end
            14'd3730 : begin out <= 64'b0010101100111011001010001111111110100101001101111010100101000000; end
            14'd3731 : begin out <= 64'b0001101011110000101010100001000100010100100101001010100011100110; end
            14'd3732 : begin out <= 64'b1010101110001010001000010001001100101001100000011010101110010111; end
            14'd3733 : begin out <= 64'b0010010011010110101010000000011100011001000011100010001111000000; end
            14'd3734 : begin out <= 64'b1010011001100111001001010100111110101000110110110010100010010100; end
            14'd3735 : begin out <= 64'b1010101110100101001010010011110100011000101000011010100100001000; end
            14'd3736 : begin out <= 64'b0010101110100101000101011011001000100100001101110010101101110100; end
            14'd3737 : begin out <= 64'b1001100110111100001010010011111010101001000011101010101001100011; end
            14'd3738 : begin out <= 64'b1010001110110000001001000011010110100101011001101010100101110010; end
            14'd3739 : begin out <= 64'b1010100101010110101010100011101010100101011100000010100000011001; end
            14'd3740 : begin out <= 64'b0010100110110010101000101101110100101100000100101010100100101011; end
            14'd3741 : begin out <= 64'b0001111110001100100111100010001100101010000110100010100000111000; end
            14'd3742 : begin out <= 64'b0010101100000110001000010110101000100111111100001010101001010100; end
            14'd3743 : begin out <= 64'b1010101111111001101000010000111010101010011100001001111111111001; end
            14'd3744 : begin out <= 64'b1010011010011110101010010010001010011010110100101010100010100011; end
            14'd3745 : begin out <= 64'b0010000010000010001010001001010100101010011110101010100000110110; end
            14'd3746 : begin out <= 64'b0010010011110101101010011001100010101011000110111010100111110111; end
            14'd3747 : begin out <= 64'b1010010101110001001010011010100100100100100100110010001011000010; end
            14'd3748 : begin out <= 64'b0010010001010111101001100001100010101011000010000010011001001101; end
            14'd3749 : begin out <= 64'b0010100000100010001010001111100100100001010101110010101000010100; end
            14'd3750 : begin out <= 64'b0010100010111110001000110011100010100111010100101010010010010100; end
            14'd3751 : begin out <= 64'b0001100110110010101000111011010010101010000111111010010011110000; end
            14'd3752 : begin out <= 64'b0010100100010000100110000001100010101001001011001010011100011011; end
            14'd3753 : begin out <= 64'b0010101100101010101000100101110000100110010101000010101010110100; end
            14'd3754 : begin out <= 64'b1010101010011111101010110011000100100101001111110010100010010011; end
            14'd3755 : begin out <= 64'b1010011011000001001001001010100100100100011110011010101000100111; end
            14'd3756 : begin out <= 64'b0010011010101000101010001000010110100100011110101010100001111001; end
            14'd3757 : begin out <= 64'b0010101111110001001010001011011110101011000100100010100001010100; end
            14'd3758 : begin out <= 64'b0010101010100010101010100011111000101001111100010010100011011010; end
            14'd3759 : begin out <= 64'b1010101010101110100111100100000000100110100000011010001001111110; end
            14'd3760 : begin out <= 64'b0010010111101000001001111101110100100101001011101010101010100100; end
            14'd3761 : begin out <= 64'b1010010111000010001001111110111010100100101101110010011100010000; end
            14'd3762 : begin out <= 64'b1010001111101111001001111010000110101011001001000010100001110101; end
            14'd3763 : begin out <= 64'b1010001101100011101001000000100010100010101001011010001100010000; end
            14'd3764 : begin out <= 64'b0001010101000110001010100111111110101001011000111010101000110100; end
            14'd3765 : begin out <= 64'b0010101000101100001001011001100110101011001100000010100110101111; end
            14'd3766 : begin out <= 64'b0010100001011110001001010100111110101001001100000010100111100101; end
            14'd3767 : begin out <= 64'b0010101000011011000111011101110010100100011001001010010010010111; end
            14'd3768 : begin out <= 64'b1001110101011010001010101001001100101000100000110010101101100100; end
            14'd3769 : begin out <= 64'b0010100100000100101001110101000100100110111011100010100100011010; end
            14'd3770 : begin out <= 64'b1010101000111111101010010000111110100101110101101010101000100010; end
            14'd3771 : begin out <= 64'b1010101100110100001000010100010110010101010111000001110001011001; end
            14'd3772 : begin out <= 64'b0010101101110101101001000110111110100000010111010010101101101100; end
            14'd3773 : begin out <= 64'b1010010101011010101010001000000100100111110011111001110110011101; end
            14'd3774 : begin out <= 64'b0010011101001110000111100111000100100100001011010001011100110010; end
            14'd3775 : begin out <= 64'b1010000001101110101001110110000000100111000000111001110000101101; end
            14'd3776 : begin out <= 64'b1001100100111011101001110000010000101011111110101010100001010110; end
            14'd3777 : begin out <= 64'b1010011011111100001010011110001010101001010000001010010100110101; end
            14'd3778 : begin out <= 64'b0010100001101100101000001010010000100101100010100010101111010110; end
            14'd3779 : begin out <= 64'b0010100110100000001010110010101110100101110110011010100001101100; end
            14'd3780 : begin out <= 64'b0010011101011100001001110000010010100111001101011010011100110010; end
            14'd3781 : begin out <= 64'b1010000111001100001010110011010000101000010011100010001110110000; end
            14'd3782 : begin out <= 64'b0001110111100111101001101010110010100100101110001010011001111100; end
            14'd3783 : begin out <= 64'b1010011100001101001010100010111010101001100110011010000100101010; end
            14'd3784 : begin out <= 64'b1010011101111101001001000101010110100010100010101010100001100000; end
            14'd3785 : begin out <= 64'b1010100100011000101010100010011000101011011001100010100101101100; end
            14'd3786 : begin out <= 64'b1010101011110000101010100110101100101011001110101010100101111000; end
            14'd3787 : begin out <= 64'b1010101101101100101010001111100000101000010110011010100110011101; end
            14'd3788 : begin out <= 64'b1001100001001111101000000000011110101001011101000010100010000110; end
            14'd3789 : begin out <= 64'b1010100101111011001010100001110110101000001100101010100100001110; end
            14'd3790 : begin out <= 64'b1010000000111100101001011010010000101010011110010010000100011110; end
            14'd3791 : begin out <= 64'b1010100001110000001010000110000010011100000011010010101001100101; end
            14'd3792 : begin out <= 64'b0010011011010100101001100011010000101011111011101010101000010000; end
            14'd3793 : begin out <= 64'b0010101011101001101010001000111010101011100011110010100111101111; end
            14'd3794 : begin out <= 64'b0010011010110010101010100001011000100001101000100010101000101101; end
            14'd3795 : begin out <= 64'b0010101101001101001001000000011110101001110011100010101010111101; end
            14'd3796 : begin out <= 64'b1010100111110110001010001110100110100011010111001010010000010110; end
            14'd3797 : begin out <= 64'b0010101101001011101000000111000000100010001010111010010011110010; end
            14'd3798 : begin out <= 64'b1010100000101010101010110011100000100010001111100010100000000010; end
            14'd3799 : begin out <= 64'b0010100100101000101010001000010100100111101111111010101100111100; end
            14'd3800 : begin out <= 64'b1010011110011111001010110000010110101000100101010010010011001110; end
            14'd3801 : begin out <= 64'b1010100010001100001011000011110010101011001010011010100100010010; end
            14'd3802 : begin out <= 64'b0010100111000111101001001111000100101000000101111010101010001000; end
            14'd3803 : begin out <= 64'b1010101100010110101010010011101000100100000101010010001100000110; end
            14'd3804 : begin out <= 64'b1010100111001001001010111101001100100110101101101010101111011000; end
            14'd3805 : begin out <= 64'b0001110111110010101001111011011000011110100110100001110001001100; end
            14'd3806 : begin out <= 64'b1001111010001011101000011000001010010111000100000010011011000010; end
            14'd3807 : begin out <= 64'b0010100010011100101000111001000010100011000111101010011001000111; end
            14'd3808 : begin out <= 64'b0010011101001000100110011111101000101011100111101010101010011011; end
            14'd3809 : begin out <= 64'b1010100111110110101010011101000100100110001010100001110011010010; end
            14'd3810 : begin out <= 64'b0001000011011100101001111111000110101011000101011001111011010111; end
            14'd3811 : begin out <= 64'b0010101101000111101010001000000000100000101100011010100011010101; end
            14'd3812 : begin out <= 64'b1010011110000101101001010011010000101011001010000010001011100001; end
            14'd3813 : begin out <= 64'b0010101100101100101010011010110000100011101010111010010010110000; end
            14'd3814 : begin out <= 64'b0010010000000010101010100011111000101010101000001010100001111000; end
            14'd3815 : begin out <= 64'b1010011110000011001010110011011110101010000111110010000111100111; end
            14'd3816 : begin out <= 64'b1001011101101101001010110100000010100110100110001010010111101110; end
            14'd3817 : begin out <= 64'b0001001001010100001001111001011110101000001101011010011101111101; end
            14'd3818 : begin out <= 64'b0010100110111010001010100110110000101011000001111010010011011110; end
            14'd3819 : begin out <= 64'b0010010010110101101001011010011110101001001000101010100101101110; end
            14'd3820 : begin out <= 64'b1010100100100100001001001101010100100101000100010010101011000111; end
            14'd3821 : begin out <= 64'b1010101001110011001010011100111010100101001001010010000000000100; end
            14'd3822 : begin out <= 64'b1010001111110011101000000011011010101000011001101010101100010001; end
            14'd3823 : begin out <= 64'b1010100000001010101001000011100110101010000001111001001111101110; end
            14'd3824 : begin out <= 64'b0001101011100000101001111001010100100011101100011001101110111011; end
            14'd3825 : begin out <= 64'b1010011110001111100111000000000010101000101011101010100011011110; end
            14'd3826 : begin out <= 64'b1001100111101000000011100100010100100100101011100010011010101011; end
            14'd3827 : begin out <= 64'b0010011110010000101010100010011000100110001000101001101111001010; end
            14'd3828 : begin out <= 64'b1010100100101001101010111101100010101000110010111010000110001101; end
            14'd3829 : begin out <= 64'b0010100010111010101010100100000110101000111100010010000101110111; end
            14'd3830 : begin out <= 64'b1010110001100100001010101011000010100011100100101010100110101011; end
            14'd3831 : begin out <= 64'b1001010001000101000110000100000100101000111011001010001001000101; end
            14'd3832 : begin out <= 64'b1010100011000100101010010101100010101011101101010010100001101001; end
            14'd3833 : begin out <= 64'b0010100111100001001001001000110000101011011111110010100101101111; end
            14'd3834 : begin out <= 64'b0010101000001010001001011001000010100010111100100010101101000111; end
            14'd3835 : begin out <= 64'b1010000001000101000110010110110110100100100111111010100100110100; end
            14'd3836 : begin out <= 64'b1001110111001000101001011011010000100100000100010010101111011110; end
            14'd3837 : begin out <= 64'b0010100000001110101001000100010110100100010101101001100101100001; end
            14'd3838 : begin out <= 64'b1010100001001101001010111111111110011110000011100010101011110101; end
            14'd3839 : begin out <= 64'b0001111110001101001010110101011100100111000100010010100111011101; end
            14'd3840 : begin out <= 64'b1010100110011110001010010000111000101000100100010010101101001101; end
            14'd3841 : begin out <= 64'b1010100111000010000110101101101000101100000001100010100001000100; end
            14'd3842 : begin out <= 64'b1010100101011011000111011010111010101011110110100010101111000010; end
            14'd3843 : begin out <= 64'b0010001010101000101010010110010100100101100101010010001010001110; end
            14'd3844 : begin out <= 64'b1010011000000001101010011100010000010100010000100010101000101101; end
            14'd3845 : begin out <= 64'b1010100111100110001001111010000010100010000001011010100110010011; end
            14'd3846 : begin out <= 64'b1010100010001010001010001101000110100000011100011001110111001111; end
            14'd3847 : begin out <= 64'b0010100011001001001010100111110000100000100100001000001001101000; end
            14'd3848 : begin out <= 64'b0010011001001100001001010000011010101001111101001010100001000101; end
            14'd3849 : begin out <= 64'b1001100100101010001010011101001000101010011010011010101100111001; end
            14'd3850 : begin out <= 64'b0010101110001011001010000101001010101000000100011010100000111100; end
            14'd3851 : begin out <= 64'b0010101011001011101010010100001100100100011011110010011110111101; end
            14'd3852 : begin out <= 64'b0010101110000000001001000100100100101001010100010010101010111101; end
            14'd3853 : begin out <= 64'b0010100101000111101001001100010010101000111100011010100010001000; end
            14'd3854 : begin out <= 64'b0010100010011110101010100001010010100100000110001010101011100010; end
            14'd3855 : begin out <= 64'b1010100111101111001010000011111110100010101110111010100101101000; end
            14'd3856 : begin out <= 64'b1010010101111110101010010111111000101001011010001010001000110101; end
            14'd3857 : begin out <= 64'b1010011110011111101000010100000000101000100011001010011000000000; end
            14'd3858 : begin out <= 64'b1010100011011100001000000010101100101001111101111010100101001101; end
            14'd3859 : begin out <= 64'b0010001011000100001010100001111010100101110100001010101101000111; end
            14'd3860 : begin out <= 64'b0010010011110100100100101011011000100011001011110010011111100101; end
            14'd3861 : begin out <= 64'b0010101010101111101010100011100000100000110011000010000101000000; end
            14'd3862 : begin out <= 64'b0010010111110100001001000011011100100101110011010010010101011000; end
            14'd3863 : begin out <= 64'b0010010111101000101010011101010100011010100000110010101100101010; end
            14'd3864 : begin out <= 64'b1010011011100001101010110010101010101010011000101010101100011111; end
            14'd3865 : begin out <= 64'b0010000110101000001001101010101000100100011011011010010011101011; end
            14'd3866 : begin out <= 64'b1010011001011011100111011001101000100001101101100010101101001000; end
            14'd3867 : begin out <= 64'b0010101001100110101010010110100000100100001001111010101010101100; end
            14'd3868 : begin out <= 64'b1010101001111010101010111000010100101011011111011010101100100001; end
            14'd3869 : begin out <= 64'b0010101110000001101010100000010100100110001000101010000010000100; end
            14'd3870 : begin out <= 64'b0010101110001001101001110000101100100110100111001010001011010110; end
            14'd3871 : begin out <= 64'b0010010110111000001010001001001110100110000100100010101001110101; end
            14'd3872 : begin out <= 64'b0010100011111001000111010110111100101010001011110010100010101100; end
            14'd3873 : begin out <= 64'b1010001001111011100110110111010100101000001111001010010111011110; end
            14'd3874 : begin out <= 64'b0010101110010110101001110010110100101100000011101010101001111101; end
            14'd3875 : begin out <= 64'b0010100000100110001000101111001010101010010101010010011100001010; end
            14'd3876 : begin out <= 64'b1010101000100100001001001110111110101000111100001010010001001000; end
            14'd3877 : begin out <= 64'b1010100011011101100111011001010000101011110010111010011011111100; end
            14'd3878 : begin out <= 64'b1010010001000001101010010001101110100100000111100010001010001001; end
            14'd3879 : begin out <= 64'b0001110110111000101010100011000100100100011110100010101110001000; end
            14'd3880 : begin out <= 64'b1001101101111111101010010011101110101011010000001010100011110001; end
            14'd3881 : begin out <= 64'b1010010100001110101001000010111100100101011001101010101011011001; end
            14'd3882 : begin out <= 64'b0010100100000011001010101110111000100001111011001010001010111100; end
            14'd3883 : begin out <= 64'b1010000011111010000111101110110110100100100101100010101100111111; end
            14'd3884 : begin out <= 64'b1010100011111110101000100011001010100011101001100001110110101101; end
            14'd3885 : begin out <= 64'b0010101111011111001010100001111010101000000101010010101001011000; end
            14'd3886 : begin out <= 64'b1010011011100001101001101001101000011110110101001010101100101110; end
            14'd3887 : begin out <= 64'b1010100001111110001000110011100110101001100100110010011010110100; end
            14'd3888 : begin out <= 64'b0010001111010101001010110101010010101000010011100010100101100110; end
            14'd3889 : begin out <= 64'b0010100110111100001010111111100010101000100011000010000111100100; end
            14'd3890 : begin out <= 64'b1010101011111101101010100100110010100011001010100010011010110001; end
            14'd3891 : begin out <= 64'b0001111000100011001001000110110010101100010001100010011001011110; end
            14'd3892 : begin out <= 64'b1010100010000101101010110111000010101100000101000010101000000011; end
            14'd3893 : begin out <= 64'b0010100110110101001010111011111000100111101101010010101101001101; end
            14'd3894 : begin out <= 64'b1010001000110010001010010000100000011010111110001010010001111110; end
            14'd3895 : begin out <= 64'b1010110000000010001010001011011000101001111100011001010111001011; end
            14'd3896 : begin out <= 64'b0010101111011010001001000100100000100010001000001010010101111010; end
            14'd3897 : begin out <= 64'b0010000100010000001010110110001100101000000010111010010111111111; end
            14'd3898 : begin out <= 64'b0010010011011001100100001111101010101000010101010010011101101111; end
            14'd3899 : begin out <= 64'b0010101011110011101000011111110000100110000011100010101011001101; end
            14'd3900 : begin out <= 64'b1010010110101101000110001101110010100101001000000010100111111010; end
            14'd3901 : begin out <= 64'b0010101110100001001010001100110000101011011110000001101000011100; end
            14'd3902 : begin out <= 64'b1010100100101000101010100100100010101000110100101010101011010101; end
            14'd3903 : begin out <= 64'b1010101110001011101000000010110110100110000011010010101111100011; end
            14'd3904 : begin out <= 64'b0010100010110010001010011000111110100111110100110000111110100011; end
            14'd3905 : begin out <= 64'b1001110110101001101011000000000110101100000010111010100000101001; end
            14'd3906 : begin out <= 64'b0001111011010101101001010010110000100110100101111010011110011010; end
            14'd3907 : begin out <= 64'b1010010110000100001010001010100000101010001101001001101011000101; end
            14'd3908 : begin out <= 64'b0010100000111101001001100010110010101001000010100010100101000110; end
            14'd3909 : begin out <= 64'b1010100001111010001000101110100010101010110110111010001110101011; end
            14'd3910 : begin out <= 64'b0010101001001000101010000110010010100110011000111010100000111100; end
            14'd3911 : begin out <= 64'b0001111010001111101001000110011000101011011110011010100001011000; end
            14'd3912 : begin out <= 64'b1010001100111100101001010101010010101001101111101010100001000010; end
            14'd3913 : begin out <= 64'b1010101001000000100110110011110000101001101111001010101101010001; end
            14'd3914 : begin out <= 64'b0010010010010101001010000001101010101010110000010010010001000101; end
            14'd3915 : begin out <= 64'b0001111010110100101001100001001110101100000011011010101101000000; end
            14'd3916 : begin out <= 64'b0001100111101111101000001111000010100111100000010010100111000000; end
            14'd3917 : begin out <= 64'b0010001011011110001001101101111000101010000110011010010010010000; end
            14'd3918 : begin out <= 64'b1001110011111001101000110000111000010000100010111010100000110101; end
            14'd3919 : begin out <= 64'b1010010111010100101000110111000000101000100110010010011011010011; end
            14'd3920 : begin out <= 64'b1010010011111000000111010110100010101011000011001010100001000110; end
            14'd3921 : begin out <= 64'b1010100011100111001000000100101100100111010000100001010100010011; end
            14'd3922 : begin out <= 64'b0010100111100010101010001110011000101010101010101000110101010010; end
            14'd3923 : begin out <= 64'b0010101011011100001010111010101000101010001010000010001011111011; end
            14'd3924 : begin out <= 64'b0010101101101110100110110111111100100001100001110010000000001101; end
            14'd3925 : begin out <= 64'b0010011000000011101001010001000100101000010101000010001111101011; end
            14'd3926 : begin out <= 64'b1010100011110100101011000000100100100110010100011010101010010010; end
            14'd3927 : begin out <= 64'b1010101011101011001010001010110100100110101010001010101100110011; end
            14'd3928 : begin out <= 64'b1010000011011011001010110110111010100111000100110001101111110111; end
            14'd3929 : begin out <= 64'b0010101000001100101001111001101000101001100011010010100000001101; end
            14'd3930 : begin out <= 64'b1010101001010110101001100000001000101100000000010001111100111111; end
            14'd3931 : begin out <= 64'b1010101110010101001010111100100010101011000000100010101011101011; end
            14'd3932 : begin out <= 64'b1010101000111110101001001101111000100110100010101010101000001100; end
            14'd3933 : begin out <= 64'b0001111100011010101010111110111010100100110001011010101110010111; end
            14'd3934 : begin out <= 64'b0010101111110011101010000100111110100000010010101010000100010001; end
            14'd3935 : begin out <= 64'b1010100000001111101010010110000100101010001001111010100011011110; end
            14'd3936 : begin out <= 64'b1001111011001110001010111110001010011100011000001001011100010100; end
            14'd3937 : begin out <= 64'b1010011001110110001001001000100010101000011101101010000010110100; end
            14'd3938 : begin out <= 64'b0010100011001110101010101100001110101011001001001001100101000101; end
            14'd3939 : begin out <= 64'b0010101111100100101010010000010010100010001000111010100101100110; end
            14'd3940 : begin out <= 64'b1010101010001001000110101010100010101010100110101010011110101110; end
            14'd3941 : begin out <= 64'b0010011000100100001001111101001100101001000011011010100111010010; end
            14'd3942 : begin out <= 64'b1010100111001111101010100111101010011110000111111010001000101111; end
            14'd3943 : begin out <= 64'b0010100010000010001010010111101000101010000110111010100101010101; end
            14'd3944 : begin out <= 64'b0010101100001101101010011110110100100010000111000010000111101000; end
            14'd3945 : begin out <= 64'b1010010011111010001001011111110100101000011010010010001100001111; end
            14'd3946 : begin out <= 64'b1010010000001101001001011001001010100011011010010010011011001011; end
            14'd3947 : begin out <= 64'b0010010111100111101001000110000010100000000000000001111000000110; end
            14'd3948 : begin out <= 64'b0010011101010110100100110100110110101001000000011010100001000101; end
            14'd3949 : begin out <= 64'b0010101000100100101010000101011100101011101110001010100001000111; end
            14'd3950 : begin out <= 64'b1010000010101010001010011010111110100000000110010010100110111010; end
            14'd3951 : begin out <= 64'b1010101001010010001010110101110110001111110000011001100110010100; end
            14'd3952 : begin out <= 64'b0010100010011001101001011110011110101010101010011010010100010001; end
            14'd3953 : begin out <= 64'b0010000000101010101001011111010010101000110100011010101100101100; end
            14'd3954 : begin out <= 64'b0010100001010011101000100110111010101001001100000010001011010011; end
            14'd3955 : begin out <= 64'b1010010101110100101000010101010010101010101010101010100110010110; end
            14'd3956 : begin out <= 64'b1001111010001010101000110000011000100101111000000010001010111001; end
            14'd3957 : begin out <= 64'b0010100001010011101010100000111100101011110010110010100010000101; end
            14'd3958 : begin out <= 64'b1010010000111011001001110001001010100100101110001010101110111001; end
            14'd3959 : begin out <= 64'b0001110011001101001010100101100110101001001001011010101001100111; end
            14'd3960 : begin out <= 64'b0001110001110110101010110011011110101000100111101010101101011011; end
            14'd3961 : begin out <= 64'b0001111101111101101000100110010110101011011111011010011001100000; end
            14'd3962 : begin out <= 64'b0010100000011111101001111011010010100001110011101010101101100100; end
            14'd3963 : begin out <= 64'b0010101101111110100111111000110100101000100000101010000011001111; end
            14'd3964 : begin out <= 64'b1010101011010111001000101101100010100100011110000010100001011011; end
            14'd3965 : begin out <= 64'b0010000011100110000110010100110100011101110100100010010000111101; end
            14'd3966 : begin out <= 64'b0010010100010001001010011001101000101011100011110010010111110010; end
            14'd3967 : begin out <= 64'b0010101100011011101010000101011000100111001001001010011110110001; end
            14'd3968 : begin out <= 64'b1010100111111010101000011001101010101011001011011010010101010010; end
            14'd3969 : begin out <= 64'b1010001010101010001001011010010100100101000100110010101001001011; end
            14'd3970 : begin out <= 64'b1010010000111000001010000110000100101000111101100010000111111110; end
            14'd3971 : begin out <= 64'b1010000101010110001010101110010110100100101011100010101010010100; end
            14'd3972 : begin out <= 64'b0010001110100011001010110100000100100100100101101001110110010000; end
            14'd3973 : begin out <= 64'b0010010100001000101010011010011100100110110111000000011000011111; end
            14'd3974 : begin out <= 64'b0010100101110111101001111110101000010101011010000010101010100100; end
            14'd3975 : begin out <= 64'b0010101100111101101001100100111100101001100101001010101111001100; end
            14'd3976 : begin out <= 64'b1010000011110011001010010010011010101000000010101010010000111001; end
            14'd3977 : begin out <= 64'b1010100011101011101001010101001000101011100100010010101011001010; end
            14'd3978 : begin out <= 64'b0010100111111000101010111000010000101011011001110010100111111000; end
            14'd3979 : begin out <= 64'b0001111101000010001001000001000100101000111001011010100011110011; end
            14'd3980 : begin out <= 64'b0010010110000111101010111100111110100010000011001010000001100111; end
            14'd3981 : begin out <= 64'b1010101010110100001010010101100100100111110101111010010001011100; end
            14'd3982 : begin out <= 64'b0010100000001010101001111000001000101010011010010010101100010011; end
            14'd3983 : begin out <= 64'b0001100110100001101010011111011010100111100001100010011001000100; end
            14'd3984 : begin out <= 64'b1010010111001011001000101111010000100100111111011010100001110110; end
            14'd3985 : begin out <= 64'b1010011110001001001010101110110000101000100110110010011110010100; end
            14'd3986 : begin out <= 64'b0010000011001001001000011101110100100110010000000010011101001001; end
            14'd3987 : begin out <= 64'b1010010111011001101010110110111010101000101110001010000100100000; end
            14'd3988 : begin out <= 64'b0010010110010111000100111111101110100101111101011010100101111100; end
            14'd3989 : begin out <= 64'b0010100111010011001010011010001000101001110110001010100100001010; end
            14'd3990 : begin out <= 64'b0001100010000011101000011001010110011101010100010010011011010000; end
            14'd3991 : begin out <= 64'b1010100100000101101001100101111010100100101001100010010100000110; end
            14'd3992 : begin out <= 64'b0010101010001111001010010110011010100000001010101010100010100000; end
            14'd3993 : begin out <= 64'b1001011000110001101001111010000000101011001010011010011010111100; end
            14'd3994 : begin out <= 64'b1010100010111010101001110011011110101010000111001010100010100000; end
            14'd3995 : begin out <= 64'b1001110111001000101010000011000010100110011001010010100010111100; end
            14'd3996 : begin out <= 64'b1010101111011111000100101110001110101010001000110010101101101010; end
            14'd3997 : begin out <= 64'b1010011001001010101010000000011010011110100100111010101111100000; end
            14'd3998 : begin out <= 64'b1010101010001110001010001101001000011001110100101010101101110010; end
            14'd3999 : begin out <= 64'b1010000011101001001000010100101110011101111100010001011100101101; end
            14'd4000 : begin out <= 64'b1010010010100111100000000011000110101010010011010001111001111010; end
            14'd4001 : begin out <= 64'b0010101100011101001010010000011110101100000010100010011101001000; end
            14'd4002 : begin out <= 64'b1010001111100001001010011001011000101001000101100010100111000111; end
            14'd4003 : begin out <= 64'b0010101010101100101010010100010010011110000011000010101001000010; end
            14'd4004 : begin out <= 64'b0001110011101000001001011011011110100011010110111001100010011010; end
            14'd4005 : begin out <= 64'b0010001101110110101001011101111100101001001101000010100001010111; end
            14'd4006 : begin out <= 64'b1010101101111110101000010100111010101010101111010001011110001000; end
            14'd4007 : begin out <= 64'b0010100111011010001001000100110100101000100100101010101100111101; end
            14'd4008 : begin out <= 64'b0001110001110011001010011001011000101001101101110010101100001001; end
            14'd4009 : begin out <= 64'b0001100111100000001010111000101110101000110011110010100100011110; end
            14'd4010 : begin out <= 64'b1010100011100110101001110111011010101000100111010010101101011110; end
            14'd4011 : begin out <= 64'b1010101000001001101010100110010010101010001000111010100011101011; end
            14'd4012 : begin out <= 64'b0010010111010101001010100100110000100100111001110010100111111000; end
            14'd4013 : begin out <= 64'b0010100001000111001000100100001110101010000010001010010000001110; end
            14'd4014 : begin out <= 64'b0010101101001100001010001100000110101010001101010010010101111011; end
            14'd4015 : begin out <= 64'b1010011110000100101010110000111010101010000000001010010111111101; end
            14'd4016 : begin out <= 64'b1010010010010100101011000000000100101010011100100010010000011011; end
            14'd4017 : begin out <= 64'b1010100110010010101001000101111100100111101100100010010001011101; end
            14'd4018 : begin out <= 64'b1010010100110001101010011111100100011111000001000010011101000101; end
            14'd4019 : begin out <= 64'b1010000101001101001010111000000100011100110010000010010011111000; end
            14'd4020 : begin out <= 64'b0010010101110001101010011011101010101011000001110010010000111011; end
            14'd4021 : begin out <= 64'b1010000110011100001010100111110000101000000110011010100010001111; end
            14'd4022 : begin out <= 64'b0010101100010011101000001001100010100000111010111010011000110011; end
            14'd4023 : begin out <= 64'b1010101100100000000110010000010110011101010111101010101000110000; end
            14'd4024 : begin out <= 64'b1010100001011101001010111000111010100010101110100010100000011001; end
            14'd4025 : begin out <= 64'b0010011101111100101000000100110010101011011100101010011010100110; end
            14'd4026 : begin out <= 64'b0010100110100010101010010010010100011001110110111010001110011011; end
            14'd4027 : begin out <= 64'b1010100101110101001001001011101100100010111111100010100011001111; end
            14'd4028 : begin out <= 64'b0010010000100100001010110011100110100100111000010010101000011110; end
            14'd4029 : begin out <= 64'b1010100100000001001010010101010100100100111110001010001110101000; end
            14'd4030 : begin out <= 64'b1010010101000111101001100111110000100000011101000010100010010111; end
            14'd4031 : begin out <= 64'b0010011110010000101000100110001000101001010000011010011011100100; end
            14'd4032 : begin out <= 64'b0010010101001011001001010101100100101011101010001010010100111110; end
            14'd4033 : begin out <= 64'b1010101110110100101001101110111110100010111101000001100011000011; end
            14'd4034 : begin out <= 64'b1010001101110110101010101101011110101010010100110010010000010101; end
            14'd4035 : begin out <= 64'b1010100011110000001010101001100010100101100010011010001100110111; end
            14'd4036 : begin out <= 64'b1010100001111111101001011100101110011110101100010010100111011100; end
            14'd4037 : begin out <= 64'b1001111010110000001001110111011010100110000011100010100111100000; end
            14'd4038 : begin out <= 64'b0010101110111001001001001111011100101001001100100010010100110011; end
            14'd4039 : begin out <= 64'b1010101011110001000101011001101100011011100101111010101001111001; end
            14'd4040 : begin out <= 64'b0010010000101111101010011110001010101011100110111001111011010000; end
            14'd4041 : begin out <= 64'b0010101011011110001010110100000100101010100011001001111100100010; end
            14'd4042 : begin out <= 64'b1010000000111101001010101101000000011011010000011010101101001001; end
            14'd4043 : begin out <= 64'b0010101011101000001001010111011000100100110111111010010110001110; end
            14'd4044 : begin out <= 64'b1010010001000101100101001000011000101100000001110010010000100011; end
            14'd4045 : begin out <= 64'b0010100000001111101010011001110110101001011011001010101100110010; end
            14'd4046 : begin out <= 64'b0001110111001010001010111110100100101010010011101010101011101100; end
            14'd4047 : begin out <= 64'b0010100111000001001010001110101000011010110110001010011101101100; end
            14'd4048 : begin out <= 64'b1010100100010100001001010110000010101011110110010010001101100011; end
            14'd4049 : begin out <= 64'b1010100000010111100111011111011000100100101101000010001010001010; end
            14'd4050 : begin out <= 64'b1001110100110001101010010111101000100011001100001010101100111100; end
            14'd4051 : begin out <= 64'b1010100000111000001010011011111000011001101001000010100110100111; end
            14'd4052 : begin out <= 64'b1010101100100001101010101001101010101000101101010010001001011000; end
            14'd4053 : begin out <= 64'b0010010001101001001010101010011010100010110001011001100101110111; end
            14'd4054 : begin out <= 64'b0010010101000100000100000100100100101010010000111010000000001110; end
            14'd4055 : begin out <= 64'b0010011111111110101001010001111100100100010011011010001111010111; end
            14'd4056 : begin out <= 64'b0010101100010011101010111001110100100001000101111010101001101000; end
            14'd4057 : begin out <= 64'b0010101110110110001001011111100010101001100100100010101100100011; end
            14'd4058 : begin out <= 64'b0001101101100111001010000111101110101010010010000010010111110111; end
            14'd4059 : begin out <= 64'b0010101111000010101001010010000110101001110100010010010001011110; end
            14'd4060 : begin out <= 64'b0010101101111110001010000010011100010101001101100010011011111110; end
            14'd4061 : begin out <= 64'b0001111001101101101010110001101000100001111100010010000100011011; end
            14'd4062 : begin out <= 64'b0010000010001110101010000101000010101011110101010010101001100010; end
            14'd4063 : begin out <= 64'b1010101011111001101010001101100110011110010111100010100010101010; end
            14'd4064 : begin out <= 64'b0010011011111011001010001000010110101010111100101010101010001110; end
            14'd4065 : begin out <= 64'b1010010011011001001010000111000110101011010111110010010010011010; end
            14'd4066 : begin out <= 64'b0010011001000110001010111100101000100100001000001010010100100010; end
            14'd4067 : begin out <= 64'b0010010111111010001010110101110100100001110111000010001110101100; end
            14'd4068 : begin out <= 64'b1010101101010011100101110110111010101000100101010010101001001111; end
            14'd4069 : begin out <= 64'b0010101111001100101010001111111100100110010011001010010110110110; end
            14'd4070 : begin out <= 64'b1010010110000101101010011101110110100000000011011010001011001111; end
            14'd4071 : begin out <= 64'b0010101011111010001010101000000000101000011101011010011000010010; end
            14'd4072 : begin out <= 64'b1010101001011101001001100101000010101010101111010010100101101101; end
            14'd4073 : begin out <= 64'b0010100110101111001000100101101100011111100111000001111010100010; end
            14'd4074 : begin out <= 64'b0010100011000010000111111101110000100000100010000010010000110110; end
            14'd4075 : begin out <= 64'b1010100001111000001001001010100000101011001000110010101110101111; end
            14'd4076 : begin out <= 64'b0010101000000011001000101111011110011111001100110001011011100101; end
            14'd4077 : begin out <= 64'b0010101010011110101010110101000100100010011111010010100101100111; end
            14'd4078 : begin out <= 64'b0010000101001110101010000101101000100101100001101010101101110001; end
            14'd4079 : begin out <= 64'b1010100110110110000110111000101010100111000111000010100000110111; end
            14'd4080 : begin out <= 64'b0010100001100010001000111111011010101000100001001010101011111111; end
            14'd4081 : begin out <= 64'b0001111100010010001001000111000010100100010000110010000010001111; end
            14'd4082 : begin out <= 64'b1010101110110011001010111011111010101011010000100010100100010011; end
            14'd4083 : begin out <= 64'b1010101010001001001010111111001000100100011101010010011100101100; end
            14'd4084 : begin out <= 64'b0010011101010110001010101001000110011110100001111010000100010100; end
            14'd4085 : begin out <= 64'b0001110101111111101010011001101100100000110110101010101111110001; end
            14'd4086 : begin out <= 64'b0010001001110001001001101010111110011001101111110010010000011111; end
            14'd4087 : begin out <= 64'b0010001001000100101010011011010000101000011001001010100101100100; end
            14'd4088 : begin out <= 64'b0010101111001010101010011000010110100101101010111010000011010011; end
            14'd4089 : begin out <= 64'b1010101110100011100111110100001010101011110000101010011100101000; end
            14'd4090 : begin out <= 64'b0010000000001100001001011001001000101001110001100010010010010110; end
            14'd4091 : begin out <= 64'b1010011010010100001001100100010000101010001000110010010000101001; end
            14'd4092 : begin out <= 64'b0010100011010011101010100010001110100110100011001010100011101011; end
            14'd4093 : begin out <= 64'b0010101100101000001010100101111100100111001111001010100111011100; end
            14'd4094 : begin out <= 64'b1001111111100010101001011101111100100100110111111010010110000011; end
            14'd4095 : begin out <= 64'b1001110001011011101010000101011100011101011001001010011010011011; end
            14'd4096 : begin out <= 64'b1010100111001100001001011011001000101001010000111010100001100011; end
            14'd4097 : begin out <= 64'b0010010101101000000111011001010000011001011110011010101100001010; end
            14'd4098 : begin out <= 64'b0010101101000101001010110111011010100101111011000010010100110110; end
            14'd4099 : begin out <= 64'b1010011100001110001010011100000010001100101110101010100000111010; end
            14'd4100 : begin out <= 64'b0010010101101100101001011010010110100101101000000010101010011001; end
            14'd4101 : begin out <= 64'b0001010110101011101000100001011100101001110110101001010001100011; end
            14'd4102 : begin out <= 64'b1001111011001001001010101100001110100001001101001010010111111110; end
            14'd4103 : begin out <= 64'b0001101111100010001010001001010110100011100101000010100000000011; end
            14'd4104 : begin out <= 64'b1010001010110010101010110110011110010100001100101001110110111101; end
            14'd4105 : begin out <= 64'b0000010110101101001001100110100100101001001111010001111110110100; end
            14'd4106 : begin out <= 64'b0010010100111010101010011111000000101000010100011010101000111000; end
            14'd4107 : begin out <= 64'b0010101000001010001010100111000100100101010011000010100101111100; end
            14'd4108 : begin out <= 64'b1010000101100100001000110100100100100111011101111010000000000010; end
            14'd4109 : begin out <= 64'b0010001001100111101010011100011110100111110111111010101010101000; end
            14'd4110 : begin out <= 64'b0010100100000000001010101111011100101000011111100010010001010010; end
            14'd4111 : begin out <= 64'b1010101100010100001001100101100010101010111110110010101111001011; end
            14'd4112 : begin out <= 64'b1010011111011001001000100101111110101010011001100010011011010001; end
            14'd4113 : begin out <= 64'b1010101111110111101010001100100010100111101110111010101101111000; end
            14'd4114 : begin out <= 64'b1010100000101000100111100100001010100000000110000010101011000000; end
            14'd4115 : begin out <= 64'b1010001101110101101010000011001100101001100110101010001111001101; end
            14'd4116 : begin out <= 64'b0010011110001011001001011100101110101001110010011010011001011010; end
            14'd4117 : begin out <= 64'b0010001011111110101010010111111000101010100111110001111011011001; end
            14'd4118 : begin out <= 64'b1010101110100000101010010110010000101011001000100010001011011100; end
            14'd4119 : begin out <= 64'b1010011101000101001010000110010110100111110010010010101110011110; end
            14'd4120 : begin out <= 64'b1010001111010001101010100100101100100000001010110010100110101110; end
            14'd4121 : begin out <= 64'b0010011001010000101010011010001000101010110001110001000000000001; end
            14'd4122 : begin out <= 64'b0010011111100000001010010010001100101001111000101010011010000010; end
            14'd4123 : begin out <= 64'b1010010110011101001010111011110000100010000011101001011110100010; end
            14'd4124 : begin out <= 64'b1010100011111101001001011111101100011010000110110010000111010001; end
            14'd4125 : begin out <= 64'b1010010100110100100110110000111010100100001110001010010000010110; end
            14'd4126 : begin out <= 64'b1010101000110111001011000001000100101000011010010010011010110000; end
            14'd4127 : begin out <= 64'b0010100000000011101000001001011100101010001001001001101101000100; end
            14'd4128 : begin out <= 64'b1010100111011101101010111010100000101000010010110010001000010100; end
            14'd4129 : begin out <= 64'b1010101011011101101010100000111000101001000011101001000101011101; end
            14'd4130 : begin out <= 64'b0001100111110000101001101110001100100111110001101010010110111101; end
            14'd4131 : begin out <= 64'b0010101001001100001011000001111100010010110100001010000010000000; end
            14'd4132 : begin out <= 64'b0010100001110101001000111100010110101000101011100010011001011001; end
            14'd4133 : begin out <= 64'b1010101001101010001010001100010110100110001100100001101001101011; end
            14'd4134 : begin out <= 64'b1010010111110011101001010011101000100110000011111010010110010111; end
            14'd4135 : begin out <= 64'b1010001110000010101010111011001010101000011100010010011011111010; end
            14'd4136 : begin out <= 64'b0010011011000101001010001001110010101000101101010010011011111011; end
            14'd4137 : begin out <= 64'b1001100101001111001010000110011010101001111101111010010101110101; end
            14'd4138 : begin out <= 64'b1010100100001010001010100111011100010010101011100001110111000110; end
            14'd4139 : begin out <= 64'b0010100101100010001010101101011010010100011010011010100110010100; end
            14'd4140 : begin out <= 64'b1010100011100011101010000000000000101000100100101010101001000111; end
            14'd4141 : begin out <= 64'b1001010111100010000100111001000110101010010110100001110110110110; end
            14'd4142 : begin out <= 64'b0010100011011100101010110001100000101000111111111010100010100110; end
            14'd4143 : begin out <= 64'b1010101001111001001000011001000000100100011000110010100011111001; end
            14'd4144 : begin out <= 64'b0010011101000001001010000001110010101000101110000010101101001011; end
            14'd4145 : begin out <= 64'b0010101001011101001010110000101110101000111000001010001100010010; end
            14'd4146 : begin out <= 64'b1010000100001001001010011100000000100101011000111010101010100001; end
            14'd4147 : begin out <= 64'b0010101011001001101010101111100110011101001101000010101000110100; end
            14'd4148 : begin out <= 64'b1010100001010011101000000001110000100011110110100010100010101110; end
            14'd4149 : begin out <= 64'b0001010010101011001000011111101110101001100011110010101100101000; end
            14'd4150 : begin out <= 64'b0010100010111111101000110001001100101001011101101010101111010000; end
            14'd4151 : begin out <= 64'b1010100110100110101010111100100100100110000100100010000010001010; end
            14'd4152 : begin out <= 64'b1010010110111000101010000010000100101000100000101001100001010010; end
            14'd4153 : begin out <= 64'b1001001111111000001010111110011100100000001101101010101111010100; end
            14'd4154 : begin out <= 64'b1010101011001110001001101110101100101010111110001010101001000000; end
            14'd4155 : begin out <= 64'b1010011001110011000111010110110110100110110110011010000011110000; end
            14'd4156 : begin out <= 64'b1001100011000010001001001110111010101001110001010010100111110001; end
            14'd4157 : begin out <= 64'b1010001011100001101010011000100100101011000101010010100011000100; end
            14'd4158 : begin out <= 64'b0010010000011101101010000110010000101000111000011010100000001100; end
            14'd4159 : begin out <= 64'b1010100111101100101000111000100110101010000000001010101101100101; end
            14'd4160 : begin out <= 64'b0001101010101110001000010011001000101010101010011010100001001010; end
            14'd4161 : begin out <= 64'b1010101110001001101010101011110000101001000101010010100000000001; end
            14'd4162 : begin out <= 64'b0010011010101110101001111110111100100100000001010010100001110001; end
            14'd4163 : begin out <= 64'b0010010111100111101010011010000100101010100000100010011001111100; end
            14'd4164 : begin out <= 64'b1010101101100001100111101101100110100001101101111010001010100111; end
            14'd4165 : begin out <= 64'b0010101001010111101010001110000100100011000100100010000101111110; end
            14'd4166 : begin out <= 64'b0010000110001011001010100110110110101000110111001010101010111101; end
            14'd4167 : begin out <= 64'b0010001101000100101000010110110000100010100000101010100111010011; end
            14'd4168 : begin out <= 64'b0010101111100001001010010111001110100000010100101010100110111101; end
            14'd4169 : begin out <= 64'b0010001010011000100111001000010110100000101111100010100110111100; end
            14'd4170 : begin out <= 64'b0010000101101100001010000001001100101010100010010010010101101111; end
            14'd4171 : begin out <= 64'b0010101011010010001001011110111000100100001000010010100111111100; end
            14'd4172 : begin out <= 64'b1001101111110110001010001101101010101001010010110010101101101100; end
            14'd4173 : begin out <= 64'b1001011000110101001010000010010000101011010010100010101000001011; end
            14'd4174 : begin out <= 64'b1010001110111111101010000011011000101010101111011010101001100110; end
            14'd4175 : begin out <= 64'b0001110100101110000111000111000110101010011110101010010111100111; end
            14'd4176 : begin out <= 64'b1010011010010110101010011110001110100000111011001010101010011110; end
            14'd4177 : begin out <= 64'b0001111101101101001000001110000110101011111010110010101010100010; end
            14'd4178 : begin out <= 64'b0010100101100101001001110000010010101000011011001010011101111000; end
            14'd4179 : begin out <= 64'b0010000111000000001010001101110000101001011010100010000001101111; end
            14'd4180 : begin out <= 64'b0010011110110100001010111100001010011110100011101010101111000000; end
            14'd4181 : begin out <= 64'b0010000100010110100111000110010010011100011111001010100111011101; end
            14'd4182 : begin out <= 64'b1010100100010011101000011010111100101010010011011010101100110001; end
            14'd4183 : begin out <= 64'b0010101101101111101001000101011110101010011000110010010101100111; end
            14'd4184 : begin out <= 64'b0010101001100111001010001111011100100100010001010010101001001011; end
            14'd4185 : begin out <= 64'b0010101110100111101001110100010110101010011001101010000111100100; end
            14'd4186 : begin out <= 64'b1010011011101101001010101110111000101000011001010010011111111110; end
            14'd4187 : begin out <= 64'b1010100110001011001010100010101110011101010100100010100010000111; end
            14'd4188 : begin out <= 64'b0001101101110111001010111000110110101001111011000010100011010010; end
            14'd4189 : begin out <= 64'b0010101011001011001001111110100010101000011000011010010011000011; end
            14'd4190 : begin out <= 64'b1010010100001111100110010011110010011001010101111010010000100101; end
            14'd4191 : begin out <= 64'b0010010100011101001010010000101100101010110110100001111001110100; end
            14'd4192 : begin out <= 64'b0010101011110110101000001000101110101011000110110010011000110010; end
            14'd4193 : begin out <= 64'b0010101010110010100011111111101110101011101110110010101110000100; end
            14'd4194 : begin out <= 64'b1010101101000111001000000011000010101000110011110010001011101100; end
            14'd4195 : begin out <= 64'b0010101011111111001010011100110010101000110101010001111000000101; end
            14'd4196 : begin out <= 64'b1010010110100101101010011010011100011001100011110010101000100011; end
            14'd4197 : begin out <= 64'b1010100010000000001001000000010010101001110001000001111101011011; end
            14'd4198 : begin out <= 64'b1010010110001101101010100001110100100111010111011010100010010101; end
            14'd4199 : begin out <= 64'b1010100110101100101001011010011110101100000101111010000100110111; end
            14'd4200 : begin out <= 64'b0010100100011011101010010100111100101000100001111010101000110111; end
            14'd4201 : begin out <= 64'b1010101011000000001000010010010000100000000001000010100110010000; end
            14'd4202 : begin out <= 64'b0010101111110101101010110011000100101010001000111010011110100111; end
            14'd4203 : begin out <= 64'b1010011101111110000110110101100110101011111011001010010111110111; end
            14'd4204 : begin out <= 64'b0010001001111100101010101111110110100111000101110010100101101100; end
            14'd4205 : begin out <= 64'b1001000110011101001010000110111000101011100001100010100011000001; end
            14'd4206 : begin out <= 64'b1010101110110100101010110111011100101010010111100010011011000011; end
            14'd4207 : begin out <= 64'b0010100110110001100110111111001110101011001100000010011010010101; end
            14'd4208 : begin out <= 64'b1010101000011010100111111100110110101001010100010010011011001000; end
            14'd4209 : begin out <= 64'b1010010100100100001010110101101110001101100000001010001111011011; end
            14'd4210 : begin out <= 64'b1010011101111110001010110001100010101000010101110010101110000100; end
            14'd4211 : begin out <= 64'b0010010001000000001001111100011010010110101011101010101111000101; end
            14'd4212 : begin out <= 64'b1010010111100101001001111111011110101000011011010010100001101001; end
            14'd4213 : begin out <= 64'b1010000011001100101010011000100110100011111010001010101011101010; end
            14'd4214 : begin out <= 64'b1010010001001000101001100000010100100110111010011010101010001111; end
            14'd4215 : begin out <= 64'b0010101011100000001001100111101100100100110100100010101001011100; end
            14'd4216 : begin out <= 64'b0010100110101100101001100101001100011100000001001001111111100110; end
            14'd4217 : begin out <= 64'b1010101111000001001000110010111100101010001111100010100010010101; end
            14'd4218 : begin out <= 64'b1010100011100011001010111001100110100100011010010001111101110010; end
            14'd4219 : begin out <= 64'b1010011101111001001010011110011100100111000010011010001010000000; end
            14'd4220 : begin out <= 64'b1010100100011010100110000111000110100110100100110010100110000101; end
            14'd4221 : begin out <= 64'b1010100010000100101000110011110100101000110111101010010101110110; end
            14'd4222 : begin out <= 64'b0010101011000101101000011001100100101010100001101010010110000111; end
            14'd4223 : begin out <= 64'b1010011100101000101000111000011100101011010100111010101001101010; end
            14'd4224 : begin out <= 64'b1010101111100111101000101100110010100101100100100010010001110111; end
            14'd4225 : begin out <= 64'b0010101101010001001010001010010010011011010110001010101010010001; end
            14'd4226 : begin out <= 64'b1010100111111011000110000110110100100101111010101010100011101101; end
            14'd4227 : begin out <= 64'b1010101001001001101010100101110100100101110101100001100011001111; end
            14'd4228 : begin out <= 64'b1010101001110001101000110011010000100010000001010010101100010010; end
            14'd4229 : begin out <= 64'b1010011000111010001001111111001010100110110111000010100001101000; end
            14'd4230 : begin out <= 64'b1001011110011001000100000111100100101010010011111010101000101001; end
            14'd4231 : begin out <= 64'b1010011100100101001001110111001110100000001110100010100010110100; end
            14'd4232 : begin out <= 64'b1010101111010100001010010010101110100101001011011010100101011110; end
            14'd4233 : begin out <= 64'b0001100111100000001001100000100110100011110011001010101011101110; end
            14'd4234 : begin out <= 64'b0010101011100110101000100011000010100111001111111010011001111000; end
            14'd4235 : begin out <= 64'b1010101011000001001010111010100000101000000111100010100110111010; end
            14'd4236 : begin out <= 64'b1010010110101001101010001101100100100110101000010010010111011011; end
            14'd4237 : begin out <= 64'b0010101001001010001000110011101000100110000000100010011110111011; end
            14'd4238 : begin out <= 64'b1010100110111010000110100100111100011100111000010010010000001000; end
            14'd4239 : begin out <= 64'b0010011111000100001010111110000100101000111110101010101110000000; end
            14'd4240 : begin out <= 64'b1010011001110011101010100001000100101000010010100010100011111011; end
            14'd4241 : begin out <= 64'b0010100000101010101001010011011110101010101110010010100000111101; end
            14'd4242 : begin out <= 64'b0010100110111010100111000011000100100100000111100010000001101000; end
            14'd4243 : begin out <= 64'b0010100000111011101001101101010100101000011101111010011010011010; end
            14'd4244 : begin out <= 64'b1010100101101010101010101000011000011001001001111010100100001101; end
            14'd4245 : begin out <= 64'b1010100011101010101000000110010110011111111000010010001100110110; end
            14'd4246 : begin out <= 64'b0010001001001111000000000100101100100101001101001010101111001110; end
            14'd4247 : begin out <= 64'b1010101110100100101011000001111000101010111111101010011100011111; end
            14'd4248 : begin out <= 64'b0010100000100111101000011111111100100001001000110010100110100101; end
            14'd4249 : begin out <= 64'b0001011010000111101000111000000000100111101011101010101010001000; end
            14'd4250 : begin out <= 64'b0010001011111000101010000101011100011011110010001010011001100010; end
            14'd4251 : begin out <= 64'b0010011111100001101010110110010000101010000010100010011000001110; end
            14'd4252 : begin out <= 64'b1010101101100110101010010100001110100100001111101010100011010010; end
            14'd4253 : begin out <= 64'b0001101001000110101010011011011000100011001010001001100001111100; end
            14'd4254 : begin out <= 64'b0010101110100001101000001000011100101010110010111010100011111111; end
            14'd4255 : begin out <= 64'b1010101111110111001001111001001000101011000101011010100010000000; end
            14'd4256 : begin out <= 64'b1010101101111100001010011110111010101000000100010010011000110011; end
            14'd4257 : begin out <= 64'b0001111011111111001010001101010110011100000011100010100100110000; end
            14'd4258 : begin out <= 64'b1010100110100011101001100001101100100111000110011010011110111000; end
            14'd4259 : begin out <= 64'b1010000011101000101010101111010000101010110010000010100111110001; end
            14'd4260 : begin out <= 64'b0010010010000011001010110011111110101001011111101010101001101101; end
            14'd4261 : begin out <= 64'b1010010011101000101010001001010000101000000001001001110000001010; end
            14'd4262 : begin out <= 64'b0010001011110110101001101010000110101010101010010010100001000101; end
            14'd4263 : begin out <= 64'b1010101001110111001010110010100110100010110000000010011000010011; end
            14'd4264 : begin out <= 64'b0010100001010110101010100100100010101001001010110010101010110100; end
            14'd4265 : begin out <= 64'b1010010001101100101010010011011010100010001000110010101100001011; end
            14'd4266 : begin out <= 64'b1010010011101110101001111110110000011001100110010001111101111011; end
            14'd4267 : begin out <= 64'b0010101110010110101010000011110100101000111011001010101100110011; end
            14'd4268 : begin out <= 64'b1010011111111110101010110111011000101010111001010010101011001011; end
            14'd4269 : begin out <= 64'b0010101101100010101010010111110100101000111011001010101100000110; end
            14'd4270 : begin out <= 64'b1010010001000111101010100110001100101000000100100010010001111000; end
            14'd4271 : begin out <= 64'b0010101101011110101010111011110110101011110110100010001011101100; end
            14'd4272 : begin out <= 64'b1010011000111010101001101110101110011100011001111010001100101011; end
            14'd4273 : begin out <= 64'b1010100100100110001010100011100010101001000010100010101111101100; end
            14'd4274 : begin out <= 64'b0010011011111111101010100111010110101010001110010010001101110000; end
            14'd4275 : begin out <= 64'b1010001001001010001010111010000110001100011001000001110100000001; end
            14'd4276 : begin out <= 64'b1001101101001100101001101011000100101001101011000010100000110011; end
            14'd4277 : begin out <= 64'b1010011101000111101010011110010110011011100010110010101100001011; end
            14'd4278 : begin out <= 64'b1010101100011011101010011000010100101000111111100010100110111010; end
            14'd4279 : begin out <= 64'b1010001110111101101010100001000000101001111101001010101011100000; end
            14'd4280 : begin out <= 64'b0010001101000001101001101110101100010101011011101001100001110000; end
            14'd4281 : begin out <= 64'b1010100000011000001010100100011100100111001100000010101101001001; end
            14'd4282 : begin out <= 64'b0010100100110001001010101000111100101001111010110010100110011101; end
            14'd4283 : begin out <= 64'b1010100000000011001010001100011110101000111010110010101100100110; end
            14'd4284 : begin out <= 64'b0010001100001011101010110111111010010110001101001010011001110111; end
            14'd4285 : begin out <= 64'b1010101000110101101010100111000010101001011001111010001010101110; end
            14'd4286 : begin out <= 64'b1001101000100011101010000111000010011100000010000010101000110111; end
            14'd4287 : begin out <= 64'b0010011110010000101001001001101000101001110110011010010011110011; end
            14'd4288 : begin out <= 64'b1010101110111010100101100101101000100011100110010010011011110000; end
            14'd4289 : begin out <= 64'b0010101100001100100110010011110010101011001110010010001111001100; end
            14'd4290 : begin out <= 64'b1001010000100011001010010111010100101001100010110010101100100101; end
            14'd4291 : begin out <= 64'b0010101010101101001010101100001110101011001011000010100010100111; end
            14'd4292 : begin out <= 64'b1010011011111101001000010001100100101011011111101010100000011001; end
            14'd4293 : begin out <= 64'b1001111101101001101010111011100010100100010001101010010111111001; end
            14'd4294 : begin out <= 64'b1010101011000110001010110010110110011111100010001010011011110011; end
            14'd4295 : begin out <= 64'b0010011010101011101010110010000010100110111000110010101011011010; end
            14'd4296 : begin out <= 64'b0010010100001001000111101100110110100101110110000010011110111010; end
            14'd4297 : begin out <= 64'b1010100110111010001010011010011100101010100110111010010011100100; end
            14'd4298 : begin out <= 64'b1010010101001111101010111001000000101011011000111010010010111011; end
            14'd4299 : begin out <= 64'b0010101010000101000101111110110000100100010000001010100010001010; end
            14'd4300 : begin out <= 64'b0010001001001101101010011111010110100001110000110010110000000101; end
            14'd4301 : begin out <= 64'b1010101110010110101010101001110100101000001011011010101000011000; end
            14'd4302 : begin out <= 64'b0010001000111010001001111000100010011111001101001010100010011011; end
            14'd4303 : begin out <= 64'b0010101000000010001010011001110100101001011110001010011100000011; end
            14'd4304 : begin out <= 64'b1010011110001011001001000100010010100010011010011010011011011100; end
            14'd4305 : begin out <= 64'b0010100011101110101010001011000110100001010001100010010010010000; end
            14'd4306 : begin out <= 64'b1010100011100000101010001000000000100100010101110010001100001111; end
            14'd4307 : begin out <= 64'b0010011010101100100111001011011000100001111111101010101101110110; end
            14'd4308 : begin out <= 64'b1001100111010111001001110100011110100101001100000010101110011111; end
            14'd4309 : begin out <= 64'b1010101001011101001001000101101010100111110001111010000110010101; end
            14'd4310 : begin out <= 64'b0010000101000011001001111011001110100110001100010010010100001010; end
            14'd4311 : begin out <= 64'b1010101101100000001010011011000100101001100100011010100110101000; end
            14'd4312 : begin out <= 64'b1010011010011110101001000100001110101011111010010010010001011101; end
            14'd4313 : begin out <= 64'b0010010011101111101010010110000000011100010110011001011000110010; end
            14'd4314 : begin out <= 64'b1010101011101101100111001100000010100101010110111010101010110110; end
            14'd4315 : begin out <= 64'b1010100110011100101000001011001110101001010011111010000101010110; end
            14'd4316 : begin out <= 64'b0010010001101001101010010000001000101000110110110010011111111100; end
            14'd4317 : begin out <= 64'b1010101011001000001000111100110110101100000011000001101111001101; end
            14'd4318 : begin out <= 64'b0010100111110100001000011011110110101011011101100010101100000101; end
            14'd4319 : begin out <= 64'b0010000011100010101001111100101000100000100010110010101000011001; end
            14'd4320 : begin out <= 64'b0010011111111010001001011110100110101001100111110010101011101011; end
            14'd4321 : begin out <= 64'b1010101010111101101001111011101010010110000100100010000011001110; end
            14'd4322 : begin out <= 64'b0010010101011000000010101100011000101100000110000010010010110111; end
            14'd4323 : begin out <= 64'b1010100100000110001010001101010000101010000000001010100110111101; end
            14'd4324 : begin out <= 64'b0010101111101000101010000101001100101010010101100010011100011000; end
            14'd4325 : begin out <= 64'b0010010001000011100110010010011100010100010101011010010100100110; end
            14'd4326 : begin out <= 64'b0010101000100011000111000011101000101010100011100010010011101000; end
            14'd4327 : begin out <= 64'b0010100010000101100011011001110000100100111101111010101011010100; end
            14'd4328 : begin out <= 64'b1010100101001001101010000000000110101000110011010010100101000111; end
            14'd4329 : begin out <= 64'b0001100001111000001010101111110010101001010110101010100001110011; end
            14'd4330 : begin out <= 64'b0001110101000000001010000100100010100110111001001010011110110011; end
            14'd4331 : begin out <= 64'b0010101001001101001010101000000000101000111001111010100010000110; end
            14'd4332 : begin out <= 64'b0010000001110010100111111111010100100001111001111001101010011111; end
            14'd4333 : begin out <= 64'b1010101000010000101010001100001010100100011101011001111110011111; end
            14'd4334 : begin out <= 64'b0010100110111000001000000101111110100110111111001010100101000000; end
            14'd4335 : begin out <= 64'b1010101011010100101010010110100000100000111011001010001011100000; end
            14'd4336 : begin out <= 64'b0010101111111101001001010111100010001101011110010010101110010001; end
            14'd4337 : begin out <= 64'b1010100110011011000111010111111110100101000000011010101011010100; end
            14'd4338 : begin out <= 64'b1010100110100110101010001001100010100111011111100001111100000010; end
            14'd4339 : begin out <= 64'b0010101110111110101000111101101100011011100101000010101010101101; end
            14'd4340 : begin out <= 64'b0010100010111010001001000101011010100000010111101010101111100010; end
            14'd4341 : begin out <= 64'b0001101100001011101010110001010000101000011110011010011010011011; end
            14'd4342 : begin out <= 64'b0010000110101111001011000000100010100001111011000010010110010100; end
            14'd4343 : begin out <= 64'b0010101100010001101000111100001100100110110100010010000011001111; end
            14'd4344 : begin out <= 64'b1010100110001000001001000001100000100011000001001010011000101011; end
            14'd4345 : begin out <= 64'b0010101110111011101010101011010100101011001000000010010010101111; end
            14'd4346 : begin out <= 64'b1010010100110001001000001111011100101001110111100010101000011001; end
            14'd4347 : begin out <= 64'b0010000110111010101010110100111100101011111010111010101110001111; end
            14'd4348 : begin out <= 64'b0010010011011000101010011110000010011111111111111010100101011100; end
            14'd4349 : begin out <= 64'b1010101010110100001001001110111110101010100111010001110111010001; end
            14'd4350 : begin out <= 64'b1010101001100010001010101100001000100010110011001010100111100110; end
            14'd4351 : begin out <= 64'b1010100010110101001010101000011000101001011010111010011011110000; end
            14'd4352 : begin out <= 64'b0010011000010101101010110101011110100100010100101010011111001110; end
            14'd4353 : begin out <= 64'b0010100101011010001001110110010000101000011101010010010011001011; end
            14'd4354 : begin out <= 64'b1010101011110010100000100011001010011101001001101010001101110011; end
            14'd4355 : begin out <= 64'b0010000101010001101010011000100010101000001101101010100011110110; end
            14'd4356 : begin out <= 64'b1010001010010000100111010101010100100111110110101010011101010110; end
            14'd4357 : begin out <= 64'b1010000110111001001000001000101010010111111011010010101111000111; end
            14'd4358 : begin out <= 64'b1010000011000010100101100110111100100000110011010010100111011110; end
            14'd4359 : begin out <= 64'b1010100010001011101010001011101100100000111011111010100010100101; end
            14'd4360 : begin out <= 64'b0010010110011011101010001001001000100101001011000010011010111100; end
            14'd4361 : begin out <= 64'b0010010111100101101010010100101110101011001100101010101101011111; end
            14'd4362 : begin out <= 64'b1001110111010010000111010100110010011101011101001010001011101010; end
            14'd4363 : begin out <= 64'b1010101011000111001010011110100000101011111010101010000111110011; end
            14'd4364 : begin out <= 64'b1010100110100100001001010111001000101010000101011010001010111110; end
            14'd4365 : begin out <= 64'b0010101100100000001000110101011100101001100011100010100101000000; end
            14'd4366 : begin out <= 64'b0010011100011000101010000011100100101000000111100010100001000111; end
            14'd4367 : begin out <= 64'b0010001010110001101001110100001000100010110010110010100110011010; end
            14'd4368 : begin out <= 64'b1010010101001011001010110001100010100110101011001010100101000011; end
            14'd4369 : begin out <= 64'b0010011000101101001010011001110000101001110111010010101100101101; end
            14'd4370 : begin out <= 64'b0010010101101000001000010001100100100000001111101001010000110001; end
            14'd4371 : begin out <= 64'b0001011010100101101001011110000100101001011010110010100011101101; end
            14'd4372 : begin out <= 64'b0010100110001010001010010110011110101001111111001010101101100011; end
            14'd4373 : begin out <= 64'b1010011110101001100111000010011100100010100110101010010001100010; end
            14'd4374 : begin out <= 64'b1010101110100100001001100101001100101001010001011010101111101100; end
            14'd4375 : begin out <= 64'b0010100111000111001010110111010000100000000110001010100000111110; end
            14'd4376 : begin out <= 64'b0010010111010101000100000110000000011101010000000010100000001011; end
            14'd4377 : begin out <= 64'b1010011011110111001010000001011100100110010011110010100100011000; end
            14'd4378 : begin out <= 64'b0010100001111000101001101000111100101011101110000010011010010000; end
            14'd4379 : begin out <= 64'b0010101110010101101010101100001110100011011001011010011001111111; end
            14'd4380 : begin out <= 64'b1010100110100111000111011011010110101010001011011010010100100000; end
            14'd4381 : begin out <= 64'b1010100101100000000011110011111100101011001110011010101010011111; end
            14'd4382 : begin out <= 64'b1010100110010001101001111010110110100110100010101001111100010100; end
            14'd4383 : begin out <= 64'b1010101101010011101010010001010010101010110011011010000101000010; end
            14'd4384 : begin out <= 64'b0001000010111011101010100001100010101010000101010010011010110010; end
            14'd4385 : begin out <= 64'b0010101100100011101010111101010100100001000001101010100100111110; end
            14'd4386 : begin out <= 64'b0010101000011101101010110010100110101000001111001010101110111100; end
            14'd4387 : begin out <= 64'b0010101111100011001010110010001110100011100101110010010011110110; end
            14'd4388 : begin out <= 64'b1010101000100010001010101010010000101000011110001010101100011110; end
            14'd4389 : begin out <= 64'b1001110111000011101010000011110010101000100100001010000001010011; end
            14'd4390 : begin out <= 64'b0001111100110010001010001111101100101001110100001010101011110010; end
            14'd4391 : begin out <= 64'b1010000000001011101010000111110000010101101011011010100000011000; end
            14'd4392 : begin out <= 64'b1010100100011000101001001110101010101010010110111010010010100011; end
            14'd4393 : begin out <= 64'b0010100010011110001010000001101000100101000111000001101011010111; end
            14'd4394 : begin out <= 64'b1010011101001011101011000001011010011111110100111010101101000000; end
            14'd4395 : begin out <= 64'b0010100111011111000011000011100000101001010010110010110000010110; end
            14'd4396 : begin out <= 64'b0010100101001001100101011010001000100101011110010001100110001001; end
            14'd4397 : begin out <= 64'b0010100100110101001001110110000110100100101000100010010001110010; end
            14'd4398 : begin out <= 64'b0001111101100000001011000001101110100110001101110010101111001011; end
            14'd4399 : begin out <= 64'b1010011001110001100100011111011110101001000110010010100010011100; end
            14'd4400 : begin out <= 64'b0001101111111010101010010010111010011110000010001010100011010101; end
            14'd4401 : begin out <= 64'b1010001110110011001001111101111100100110111010101010101000111111; end
            14'd4402 : begin out <= 64'b1010101101001110001000001110000110101001010100011010011010001010; end
            14'd4403 : begin out <= 64'b0000111000111001101001000010000010100001100001000010010101010110; end
            14'd4404 : begin out <= 64'b0010010011101111101010000100101000011111100011011010100000110110; end
            14'd4405 : begin out <= 64'b0010010101110110001010110111010100011111000011110010101110111110; end
            14'd4406 : begin out <= 64'b0010101001110110101000000011111110101011111101001010101110111111; end
            14'd4407 : begin out <= 64'b1001101101100101001010100010101100100010100100010001110011101100; end
            14'd4408 : begin out <= 64'b0010010001011000101010110011001000100010110100110010101011101111; end
            14'd4409 : begin out <= 64'b0010100000101100001001110100101100101000111100110010100101110100; end
            14'd4410 : begin out <= 64'b1010100110001100101010110101011110101000000001101010100001110111; end
            14'd4411 : begin out <= 64'b0010101110000111100111111001000010100111001111101010101001111110; end
            14'd4412 : begin out <= 64'b1010100101011010101010100000110100100101101000101010101110000110; end
            14'd4413 : begin out <= 64'b0010010000100011101001010001110110100001010010101010000111000111; end
            14'd4414 : begin out <= 64'b0010100001001000101000101001110100011110011001100010100001000010; end
            14'd4415 : begin out <= 64'b0010101110010000101001100000111110101001010010001010010111100011; end
            14'd4416 : begin out <= 64'b0010100000111010001010110010101010101000001011110010101111100100; end
            14'd4417 : begin out <= 64'b0010000110001000101001101111100010101000110000000010101011010101; end
            14'd4418 : begin out <= 64'b1010101010011001000100011111110110100110000000011010100110011100; end
            14'd4419 : begin out <= 64'b0010010101001111001010001110100010100101010100000010011011000001; end
            14'd4420 : begin out <= 64'b1001110010000101001010010101110000011110001010001010101010001110; end
            14'd4421 : begin out <= 64'b1010101101100001001010110111000100100100000100101010100011001000; end
            14'd4422 : begin out <= 64'b0010000111100011100111000000011010101001001000101001111000010100; end
            14'd4423 : begin out <= 64'b1010100111010010001000100000101000101000100100000010100011000111; end
            14'd4424 : begin out <= 64'b1010101010010011101001000000110010100101111001001010100011000001; end
            14'd4425 : begin out <= 64'b0001111000011010100111111111000110101010101110101010101111000001; end
            14'd4426 : begin out <= 64'b0010100001101110001001001011110000100010011010010010100000100110; end
            14'd4427 : begin out <= 64'b1001111111111110001001100110011000101001100011101010011101100010; end
            14'd4428 : begin out <= 64'b1001100010111111001010101110110110100100011001000010000001101011; end
            14'd4429 : begin out <= 64'b0010100010110001001010010101011110101010000000111010100001110011; end
            14'd4430 : begin out <= 64'b1010010010110001001001110001010010101100001001001010101000100111; end
            14'd4431 : begin out <= 64'b0010011101110101101001100000000000101001111100110001111011000101; end
            14'd4432 : begin out <= 64'b0010010000001000101010000000101100101001111111010010000010110111; end
            14'd4433 : begin out <= 64'b1001110011000101101001101011100100101001011111000010100011001001; end
            14'd4434 : begin out <= 64'b1010011001011110001000010111111110011100001001011010101111111010; end
            14'd4435 : begin out <= 64'b1010011101000101100110111011101110101010100011100010010010011001; end
            14'd4436 : begin out <= 64'b0010000110010001101000000110001000101010101011110010100010100111; end
            14'd4437 : begin out <= 64'b1001111100001010001010101111101110100111000000001010101000000111; end
            14'd4438 : begin out <= 64'b0010011101101000101001001110011100100110001101111010000101000000; end
            14'd4439 : begin out <= 64'b1001100000111001101010110000110010100110101001010001101101110011; end
            14'd4440 : begin out <= 64'b1010001101111001101010101111110100011011011010000010010110100111; end
            14'd4441 : begin out <= 64'b0001100110101100101001101110010100100110110011001010010001111110; end
            14'd4442 : begin out <= 64'b0010101100111110001010000110000010101001111110111010011101001001; end
            14'd4443 : begin out <= 64'b1010100101011100101001000101000100101001000011101010101000101000; end
            14'd4444 : begin out <= 64'b1010100000001001000101010111101000100001010000001001111110110100; end
            14'd4445 : begin out <= 64'b0010100010110101101010101101011000101001011000010010100100110000; end
            14'd4446 : begin out <= 64'b0010010001101101101000011110010100100100101011001010011011001001; end
            14'd4447 : begin out <= 64'b0010100010110101001010101000001010101100000101101010101110010010; end
            14'd4448 : begin out <= 64'b0010100011000111000111101010100110101011000111111010100000101100; end
            14'd4449 : begin out <= 64'b0001010111001000001001011110110000100100000001110010101101110100; end
            14'd4450 : begin out <= 64'b1010100110011010101010010110001000101011001110001001110110010000; end
            14'd4451 : begin out <= 64'b1010010001011100001001010001010000101000001000001010100101001000; end
            14'd4452 : begin out <= 64'b0010101101111010001000010101101010101011101100111010011010101011; end
            14'd4453 : begin out <= 64'b0010100011011010101010001101011000101000110111011010101010101011; end
            14'd4454 : begin out <= 64'b0010010001110100101010110000111000100101010011010010011111100110; end
            14'd4455 : begin out <= 64'b1010001001001011001000101011100110101001110100011010100011100100; end
            14'd4456 : begin out <= 64'b0010101110110011101010101011101010100010111100000010101000110011; end
            14'd4457 : begin out <= 64'b1010011101110110100101101010010000101000011110100010101010100001; end
            14'd4458 : begin out <= 64'b0010100010110101100110001100010000101010110000010001110011001101; end
            14'd4459 : begin out <= 64'b1010101011011110001001010001010010100000011100010010001100010111; end
            14'd4460 : begin out <= 64'b1001110110111011001010001110000110101011010110101010011010100110; end
            14'd4461 : begin out <= 64'b0010000000111001101010101111111110100011011000110010011001111101; end
            14'd4462 : begin out <= 64'b1010100111000111001000011001010100101011111110100010100010100001; end
            14'd4463 : begin out <= 64'b1001110110111000101010010000111010101010110011101010101101100110; end
            14'd4464 : begin out <= 64'b0001110100010100001000001010100010101010110111000010100110110011; end
            14'd4465 : begin out <= 64'b0010101000111111101001100010110000101001100101011010011111110100; end
            14'd4466 : begin out <= 64'b1010100000111000101001110101010110101010001011111010101100100011; end
            14'd4467 : begin out <= 64'b0010100100111111001011000000111010100101011111010010001100100100; end
            14'd4468 : begin out <= 64'b1010010010001000001001001101111000101000101101010010100000010011; end
            14'd4469 : begin out <= 64'b0010101010110011001001000111010100101001000100100010101100101010; end
            14'd4470 : begin out <= 64'b1010101101000010001010001110001000101010011010011010101110011011; end
            14'd4471 : begin out <= 64'b0010010110110000101001000010001110101010010010001010100010111000; end
            14'd4472 : begin out <= 64'b1001110001100100101010111100011110101011111011101001101011100010; end
            14'd4473 : begin out <= 64'b0010100110000100000111001100111110100011111110010001110010100001; end
            14'd4474 : begin out <= 64'b0010101011101111101000111000100000100001101011110010000001101010; end
            14'd4475 : begin out <= 64'b0010100111111011101010001001100000101001100010011010101011111101; end
            14'd4476 : begin out <= 64'b1010011001111011001010010001100110011111101011110010011001111100; end
            14'd4477 : begin out <= 64'b1010000010010001001010011111010110101011100111001010001011001000; end
            14'd4478 : begin out <= 64'b0010100101101000101001100101011100101000000000100010010100011110; end
            14'd4479 : begin out <= 64'b0010101100011011101001000111001000011110011101101010100001111101; end
            14'd4480 : begin out <= 64'b0010101111001000001001010010101010100100010001001010011010111010; end
            14'd4481 : begin out <= 64'b1010100001111110001001000100011000100100110111100001110110000010; end
            14'd4482 : begin out <= 64'b1001100001010101001010010000010110100101010010110001110011001001; end
            14'd4483 : begin out <= 64'b1010100000101000100101101100111110100111111011111010100111110010; end
            14'd4484 : begin out <= 64'b0010101001100010101010111100100110010110101010100010101000110110; end
            14'd4485 : begin out <= 64'b0010100100110010101000100101100100101010011101100010110000001010; end
            14'd4486 : begin out <= 64'b1010100111110111001001100011100000101000100101000010101010011011; end
            14'd4487 : begin out <= 64'b1010001110100100100111011110111010000010100000010010101110010001; end
            14'd4488 : begin out <= 64'b0001111010110110000111101011110100101011010110011010100010011000; end
            14'd4489 : begin out <= 64'b1010100000000011001010000100101010100000000111000010101100010110; end
            14'd4490 : begin out <= 64'b0010011100001000000111000011010000101000101110110010000110010000; end
            14'd4491 : begin out <= 64'b0001001110101011101010110000101100101000010110011010010010110010; end
            14'd4492 : begin out <= 64'b0010101001110010101010111010100010101011111011110010101010001111; end
            14'd4493 : begin out <= 64'b1010101010100100001000100010000000011101101101010010100011110010; end
            14'd4494 : begin out <= 64'b1010101001111110101001011010110100101000001000100010101000000110; end
            14'd4495 : begin out <= 64'b0010100010000011100011110110000100011101100100010010101110111110; end
            14'd4496 : begin out <= 64'b1001101101001100000111011010010010101001010111111010011100110010; end
            14'd4497 : begin out <= 64'b0001101111010000001010110001100000101010111110110010010110111001; end
            14'd4498 : begin out <= 64'b1010100101111100101010011110010000101000010101101010001011000101; end
            14'd4499 : begin out <= 64'b0001111001010010001010010101000100100110100001110010101110110000; end
            14'd4500 : begin out <= 64'b1010100101011010001010011110101100100110100110110010100000101000; end
            14'd4501 : begin out <= 64'b1010010101111101001010000010001010100001101010111010000011110110; end
            14'd4502 : begin out <= 64'b1010001100001110101010001000101110011101011101011010011001011110; end
            14'd4503 : begin out <= 64'b0010101100110110001001110010101100100111010111101001111001001111; end
            14'd4504 : begin out <= 64'b0001100010000111101001011101101110101001100001000010010110100110; end
            14'd4505 : begin out <= 64'b0010100110101001001010111001000100101011010100110010101100101010; end
            14'd4506 : begin out <= 64'b0000111010111000100110001010000100101011110110010010000001100110; end
            14'd4507 : begin out <= 64'b1001100010011101001000111001100110100101110010101010100000110101; end
            14'd4508 : begin out <= 64'b1001111111111100001001000111101110101000101100010010010111010101; end
            14'd4509 : begin out <= 64'b1010100010000111001001000000010000100101010001010010011101100000; end
            14'd4510 : begin out <= 64'b1010011010110100001010110101111100101011011010110001010100111111; end
            14'd4511 : begin out <= 64'b0010101010100000101010001011001110100010110011101010100010101010; end
            14'd4512 : begin out <= 64'b1010101011000011101010001000111110010100100100001010010011110110; end
            14'd4513 : begin out <= 64'b1010101110001111001010000101001100100110010100100010101111001110; end
            14'd4514 : begin out <= 64'b1010001110001100001010010001111110100111101110100010011011111101; end
            14'd4515 : begin out <= 64'b1010100101101011000111111100011110101010011011110001100110010100; end
            14'd4516 : begin out <= 64'b0001110111001111101000011000111110101011100110110010100101101001; end
            14'd4517 : begin out <= 64'b0010011110100011100011001001011000100110001100111010000111110110; end
            14'd4518 : begin out <= 64'b0001111011101010000110100011000110101000100101001010010010110010; end
            14'd4519 : begin out <= 64'b0010100101010100001001100100000100100101111100111010001001000011; end
            14'd4520 : begin out <= 64'b1010011100001111101010000100110110100001110101010010100011110100; end
            14'd4521 : begin out <= 64'b0010101000000010101000100010101010100100100001101010010101011010; end
            14'd4522 : begin out <= 64'b0001101000111101000111101111010110101001011010110010000010000111; end
            14'd4523 : begin out <= 64'b1010100110100000001000101100010110100110001000001010100111010001; end
            14'd4524 : begin out <= 64'b0010010100100000101010010011000100101001010010100010010101101110; end
            14'd4525 : begin out <= 64'b1010101110000010001001101010011010101001101110101010100000110000; end
            14'd4526 : begin out <= 64'b1010100111011010001011000011100100100000000000011001111000000000; end
            14'd4527 : begin out <= 64'b0010100101010100101010010011111010101011101100110010101010111011; end
            14'd4528 : begin out <= 64'b1001011001101011100111001001101100101001100110110010011001000110; end
            14'd4529 : begin out <= 64'b1010010100110100001010000011000110101011100110001010011011110110; end
            14'd4530 : begin out <= 64'b0010000101000010101000101110110010100000001100101010101011100000; end
            14'd4531 : begin out <= 64'b0010001010001111001001111111000010101011111100001010010101111000; end
            14'd4532 : begin out <= 64'b1010010110111110101001001000000100100111000000010010100100010000; end
            14'd4533 : begin out <= 64'b0010100010100010001000101111101000101001101001111001110010010001; end
            14'd4534 : begin out <= 64'b1010011011110011100111110011110010101011110011110010100111111010; end
            14'd4535 : begin out <= 64'b0010100101110000101010001001101100100110110011010010101101111110; end
            14'd4536 : begin out <= 64'b0010010011001000101011000100011010101000110111010010011100000001; end
            14'd4537 : begin out <= 64'b1010010110010011100010110011101110101000100111001010101111000110; end
            14'd4538 : begin out <= 64'b0010101001100110101010000101010010101000111011100010000010101110; end
            14'd4539 : begin out <= 64'b1010011000011100001010000001000000101100001101001010100011100101; end
            14'd4540 : begin out <= 64'b1010100000101101001000011100011110011100000011111010011001101110; end
            14'd4541 : begin out <= 64'b0010001001101110100111100111001110101001001000101010011111100110; end
            14'd4542 : begin out <= 64'b1001010110011110101000001110101010101010100100010010101001010101; end
            14'd4543 : begin out <= 64'b1010101011010110001010110100010000101000101001011001100010000010; end
            14'd4544 : begin out <= 64'b0010101111111110001010011011111000101011110000011001100001111111; end
            14'd4545 : begin out <= 64'b0010100011110110001010011111001010100000110001001010010001011011; end
            14'd4546 : begin out <= 64'b1010000000101111101010000101100000100101110011011010011011001010; end
            14'd4547 : begin out <= 64'b1010101001110100001001111010101000100111101110111010101101110111; end
            14'd4548 : begin out <= 64'b0010100010101010101010010110010010100100000111011010101011101101; end
            14'd4549 : begin out <= 64'b1010100100001110100111110010100000100110111100011010110000010000; end
            14'd4550 : begin out <= 64'b0010000111000110101010110001111000101010000111001010011001010100; end
            14'd4551 : begin out <= 64'b1000111101010100101010001111000110101001000111010010100100010100; end
            14'd4552 : begin out <= 64'b0010100011000111101001101010010100100100011111010010100001011010; end
            14'd4553 : begin out <= 64'b0010010111011010101000101010001000101001111100010010101000010110; end
            14'd4554 : begin out <= 64'b1010010101100001001010010011001110100010101001110001100000000001; end
            14'd4555 : begin out <= 64'b1010101001101100101010011011001110101010000110011010011110111111; end
            14'd4556 : begin out <= 64'b1010101001010101001010001011010110100011110001001001110011100100; end
            14'd4557 : begin out <= 64'b0010100100011101101001110101100010100001000010011010001001101011; end
            14'd4558 : begin out <= 64'b0010011101010110001001101110010100100001010110101000101100100100; end
            14'd4559 : begin out <= 64'b0010011010100000001001100010100000101000101101100010000100011100; end
            14'd4560 : begin out <= 64'b1010100010110110001000101000001110101001000100000010000010001111; end
            14'd4561 : begin out <= 64'b0010100011010010101001100001110000101100000110010010011000101000; end
            14'd4562 : begin out <= 64'b1001110000101011101000111101110100100101110000110010100010010011; end
            14'd4563 : begin out <= 64'b1001011010100100001010000000000100100101110111010010011100110001; end
            14'd4564 : begin out <= 64'b1010101000100011101010011000100000101010101001100010101001001001; end
            14'd4565 : begin out <= 64'b0001100101111100101000001110010110101001111110101010100000110100; end
            14'd4566 : begin out <= 64'b0010011110110011001010111100010100101010111100101010100001011101; end
            14'd4567 : begin out <= 64'b0010101100001000001010001101010000100010011111111001111000000011; end
            14'd4568 : begin out <= 64'b1010100111001110101010101000101110100011111101000010010110100101; end
            14'd4569 : begin out <= 64'b1010100010101010101001100100101110100001000011101010010100001001; end
            14'd4570 : begin out <= 64'b1010010000011000000010001110000000100101100001111010011011110010; end
            14'd4571 : begin out <= 64'b0010011010000011001010001001110110100110010011100010010000110101; end
            14'd4572 : begin out <= 64'b1010101011101110101001100011010110100010010111111001011111110100; end
            14'd4573 : begin out <= 64'b0010011011010000001001011101001000101001011001100010000101101101; end
            14'd4574 : begin out <= 64'b0010000001011001101010001011100000011101110011100010100110100001; end
            14'd4575 : begin out <= 64'b1001101011010011101010110110100000101001101111111001111001100001; end
            14'd4576 : begin out <= 64'b0010010010010010001010011110101000100100011111010010100000100110; end
            14'd4577 : begin out <= 64'b1010101111010000101010011000011110101000010100011010100010100000; end
            14'd4578 : begin out <= 64'b0010100111001110001010010000100100101010000010100001101111011010; end
            14'd4579 : begin out <= 64'b0010100001011101000111110110010110100010110011010010011001100110; end
            14'd4580 : begin out <= 64'b1010100000011101101000110111101100011100100100111001111101000011; end
            14'd4581 : begin out <= 64'b0010100111010001101010001110010100101001110101001010101110101011; end
            14'd4582 : begin out <= 64'b1010101001100101101001010110001110101000010000001010100110101110; end
            14'd4583 : begin out <= 64'b0010100110100010101001010101110110100111101011011001111101111100; end
            14'd4584 : begin out <= 64'b1010100110101010001000100100101000011101000010110010010101001110; end
            14'd4585 : begin out <= 64'b1010011110100011101010011011100100101011110000010010011000001100; end
            14'd4586 : begin out <= 64'b1010100101001010001010111101001100100101001101011010010110101100; end
            14'd4587 : begin out <= 64'b1010101000000000001010101010100100101000110101110001000100101000; end
            14'd4588 : begin out <= 64'b0010101011011011101001101001110100101000001010111001001011101100; end
            14'd4589 : begin out <= 64'b1010100010000001001010110110100010100111001000110010011010011010; end
            14'd4590 : begin out <= 64'b0010000100100111001000011011011010101000001110101001111100111110; end
            14'd4591 : begin out <= 64'b0001111101000100001001100111101000101011001111010010000010100000; end
            14'd4592 : begin out <= 64'b0010000001110100001010010000100010101010100111110010101010000111; end
            14'd4593 : begin out <= 64'b0010011000001000101001101100010100100111101000001010101001110111; end
            14'd4594 : begin out <= 64'b0001111000101110101001000010000010101011110110000010010011000011; end
            14'd4595 : begin out <= 64'b1010010001111101101001111111111010101011100001110010011111111000; end
            14'd4596 : begin out <= 64'b0010001100010010101010000110111000101011000100010010100011100111; end
            14'd4597 : begin out <= 64'b1010010000000001001010010011001010101010111111101010010101100000; end
            14'd4598 : begin out <= 64'b0010010110010011001010000001010000100101010001101010101100110000; end
            14'd4599 : begin out <= 64'b1010100101010010001010001000001000100100101011111001110100111010; end
            14'd4600 : begin out <= 64'b0001110110000000001010100110011100101011111111101010011110111001; end
            14'd4601 : begin out <= 64'b1010101111101001001010010110100100101010011100000010010010101001; end
            14'd4602 : begin out <= 64'b0010101100001011101011000000011000101000000011011001111010111110; end
            14'd4603 : begin out <= 64'b0010000100111101101000111000100100101011010111111010101000010101; end
            14'd4604 : begin out <= 64'b1010010011001101101011000001111000101011001110110010011100000000; end
            14'd4605 : begin out <= 64'b1010101101101110001010110100001000100010001010101010100011110100; end
            14'd4606 : begin out <= 64'b0001111100000011000101111101010010101001011100010010101001010110; end
            14'd4607 : begin out <= 64'b1010100111010110101001000011011110101000001100000010100010010100; end
            14'd4608 : begin out <= 64'b1010000001000000001010101110011110101000111110011010101101001010; end
            14'd4609 : begin out <= 64'b0010011110110010001001101111001100100100110010100010101111011110; end
            14'd4610 : begin out <= 64'b0010101011100001101000010110010010011111101000011010101000001101; end
            14'd4611 : begin out <= 64'b1010100100111011001001000010011100100111011110110001100110010011; end
            14'd4612 : begin out <= 64'b0010101010010001100111000010110100100100111110001001111011010100; end
            14'd4613 : begin out <= 64'b0001111100100110001010010001010000101001101000101010101001010011; end
            14'd4614 : begin out <= 64'b0010100101100011101000001000011010100111001010011010000010111101; end
            14'd4615 : begin out <= 64'b0010011011101100101001101010011010101010101010001010100111010011; end
            14'd4616 : begin out <= 64'b1010011011001010001000100011000000100110110011100010101101110110; end
            14'd4617 : begin out <= 64'b0010101110101000001010011000101100100100001101000010000011101010; end
            14'd4618 : begin out <= 64'b0001110001111100001000101011111100100110011000000010001001011111; end
            14'd4619 : begin out <= 64'b0001100101100101001010100001101110101011101100110010101101010011; end
            14'd4620 : begin out <= 64'b0010011101100001001010000000111000100111110010000010101011001010; end
            14'd4621 : begin out <= 64'b1010100101101000000111110001000010101010110111011001101111000010; end
            14'd4622 : begin out <= 64'b0010001010010111100110111011000100101010010111101010001011001010; end
            14'd4623 : begin out <= 64'b1010101010001000101001110001011110101010001110111010100110100000; end
            14'd4624 : begin out <= 64'b0001111011010100101010101010110010100100111001111010011111010001; end
            14'd4625 : begin out <= 64'b1010100110111110001010100100100110101001011110011010101001001110; end
            14'd4626 : begin out <= 64'b1001110001110110101001111010110010100111100011101001110010110111; end
            14'd4627 : begin out <= 64'b1010010101010110101000001101101010100110001110111010101011110110; end
            14'd4628 : begin out <= 64'b1010001101100111000110111001111010100111110100001001000100010110; end
            14'd4629 : begin out <= 64'b0010100100000001001010101100011000101000100010010001011001100110; end
            14'd4630 : begin out <= 64'b1001111010110101101001111011101010101010110110001010101001101000; end
            14'd4631 : begin out <= 64'b1001000110111110001001000110110100010001001011010010100101010110; end
            14'd4632 : begin out <= 64'b1010101101001010101010101000001100100011111101001010100001110101; end
            14'd4633 : begin out <= 64'b0010011000010100000111101000110100100101101100100010101001001100; end
            14'd4634 : begin out <= 64'b0010101011001011001001110110110100101001111010000010101110100111; end
            14'd4635 : begin out <= 64'b1010000110010001101001000111000010100111110001101001010110110110; end
            14'd4636 : begin out <= 64'b1010101100100000000111001000100100010110110010111010101011101011; end
            14'd4637 : begin out <= 64'b1010000001011001001010011100011010100111000000111010011001110110; end
            14'd4638 : begin out <= 64'b0010101111011111001010100001100100101011000100010010101100110110; end
            14'd4639 : begin out <= 64'b1010110000000000001010011110000010101010001100010010100110000100; end
            14'd4640 : begin out <= 64'b1010010111101110000111111110000000011110111100110010001011101001; end
            14'd4641 : begin out <= 64'b1010100101000101101001000100111010101000010110100001100000101000; end
            14'd4642 : begin out <= 64'b0010010111110111001010011101001100101011010011001010100001111101; end
            14'd4643 : begin out <= 64'b0010100111111011001001000100110010100100000011010010010111001101; end
            14'd4644 : begin out <= 64'b1010000111010101101010101110010010100100100100001001010011101101; end
            14'd4645 : begin out <= 64'b0001010111101011001010110111010000100100111110001010010101011010; end
            14'd4646 : begin out <= 64'b0010100110101001101010011110110000101000110000011010011100001100; end
            14'd4647 : begin out <= 64'b0010011000000001000111101000001100101010101100001010100111000110; end
            14'd4648 : begin out <= 64'b1001100011100100101001101111101110011100000111001010100101100111; end
            14'd4649 : begin out <= 64'b1010101000000011101010011101101010101001100011110010001010101000; end
            14'd4650 : begin out <= 64'b0010001000001010101001001110000110101001110111110010011111110110; end
            14'd4651 : begin out <= 64'b1001110111011101100011100000010000100011011001000010010101111110; end
            14'd4652 : begin out <= 64'b0010100000111000001010110110001110100010110001011010101010000011; end
            14'd4653 : begin out <= 64'b0001101111000000101001101111110000101010110001110010100111000110; end
            14'd4654 : begin out <= 64'b0010100000111101001010010100101110100001111110011010101001111000; end
            14'd4655 : begin out <= 64'b0010100001100111101010100100100110101001100110000010101011000111; end
            14'd4656 : begin out <= 64'b0010011011100010001010001011100110101000001000010010001000001101; end
            14'd4657 : begin out <= 64'b1010101011001010101001110111001000100110110101101010101000011110; end
            14'd4658 : begin out <= 64'b0010101100001001001010100110010110101000110000000001000110101101; end
            14'd4659 : begin out <= 64'b0010100111111011001010001010100100101001011010000001111110010100; end
            14'd4660 : begin out <= 64'b1010001010101001101010101011011110101000100000111010101100110000; end
            14'd4661 : begin out <= 64'b0001111001011010101010000111111010011110100110100010000010001000; end
            14'd4662 : begin out <= 64'b1010100000101100001010111101011110101000101100010010101001001000; end
            14'd4663 : begin out <= 64'b1010100000010000101001011000001010100100001100101010101000010011; end
            14'd4664 : begin out <= 64'b1001110001000001001001111110010100101001011001001010100100110100; end
            14'd4665 : begin out <= 64'b1010100001101011101000000101011100100000101100101010001010000001; end
            14'd4666 : begin out <= 64'b0010101010111001001000011111111000101010110101010010101101001100; end
            14'd4667 : begin out <= 64'b1010100001000101000111000100001010101000110001100010101001011000; end
            14'd4668 : begin out <= 64'b0010100110011101101000000110010010011111011100011001101101101001; end
            14'd4669 : begin out <= 64'b1010100101110000000110001000111010011110011100001010000101001110; end
            14'd4670 : begin out <= 64'b0010101111100111101010000011011110101011011110110010100101101001; end
            14'd4671 : begin out <= 64'b0010101101110110001001101100100000100100000101010010001101011111; end
            14'd4672 : begin out <= 64'b0010000110101110101001101001001100100111010101000010101000000010; end
            14'd4673 : begin out <= 64'b0010000011001101101010000010001010101010111001000010100011000000; end
            14'd4674 : begin out <= 64'b0010101110100111001010010110010100100010001011010010100000100000; end
            14'd4675 : begin out <= 64'b1010011011111001101010101100101110101010000101000010011111101001; end
            14'd4676 : begin out <= 64'b0010001111010111001010111001111000101011001110001010011101111011; end
            14'd4677 : begin out <= 64'b0010101011011011000111001100101000100001101010010010000101110111; end
            14'd4678 : begin out <= 64'b0010100000111111001000111111001100101011000100100010001010011001; end
            14'd4679 : begin out <= 64'b0010101101100001101000011101010010011001011101000010011010110010; end
            14'd4680 : begin out <= 64'b0010100011100000001001101010101010100001001101001010101110110010; end
            14'd4681 : begin out <= 64'b1001110001110101101010000000001110101011011111100001000000001101; end
            14'd4682 : begin out <= 64'b1010011011000111101010100010110010100100111001111010011010100001; end
            14'd4683 : begin out <= 64'b1010100111001000100101010111111100101000111011111010010011100111; end
            14'd4684 : begin out <= 64'b0010100100010000000111100011111000101010001001001010000000111011; end
            14'd4685 : begin out <= 64'b1010011011001100101001110001100100100000111110100001111110110100; end
            14'd4686 : begin out <= 64'b1010101111100101101010111110000000100111100100110001100110110110; end
            14'd4687 : begin out <= 64'b0010101011000111101001000011110010100001000100111010100001010010; end
            14'd4688 : begin out <= 64'b0010101001100110001010010111110000100010011100101010100000100111; end
            14'd4689 : begin out <= 64'b1010011001010001100110011111100110100011100011000010010111100010; end
            14'd4690 : begin out <= 64'b1010000000000011001010100101010110011011011001111010100011001001; end
            14'd4691 : begin out <= 64'b0000100100010111101010101111010110101010000010100001110100110010; end
            14'd4692 : begin out <= 64'b1010011000111011000110010111000000101000001000111001101010010110; end
            14'd4693 : begin out <= 64'b0010101000111010001010011011000000101001110110101010000011101010; end
            14'd4694 : begin out <= 64'b1001111110110000001010101001111010101000111000000010100111110010; end
            14'd4695 : begin out <= 64'b1001101011110101000111101101100010100100001110000010000000100111; end
            14'd4696 : begin out <= 64'b1010010101010010001010001111011100101010001100100010010100111100; end
            14'd4697 : begin out <= 64'b0010000010000101101010011100001110100100000001000010101100110001; end
            14'd4698 : begin out <= 64'b0010001100110110001010101001000110011110001111100001100111000000; end
            14'd4699 : begin out <= 64'b1010100011111100101010000010111000100010000110111010100101011101; end
            14'd4700 : begin out <= 64'b0010110000111000101010110010000000101000111001001010011010111101; end
            14'd4701 : begin out <= 64'b0010011101101000101010111110000000101011101001110010101111101100; end
            14'd4702 : begin out <= 64'b0010000100000001101010110011010000101010001000000010100011011110; end
            14'd4703 : begin out <= 64'b0010100001100011001010100000001100101001001001110010001101011111; end
            14'd4704 : begin out <= 64'b1010101000100101001001010010010000100011111001111010100011010100; end
            14'd4705 : begin out <= 64'b0010100011010001101010000100000000100111000000000010100000111000; end
            14'd4706 : begin out <= 64'b0010010111010000001001011110000000100110011000010010100110000000; end
            14'd4707 : begin out <= 64'b1010101001110100001010100110111100101011001100100010000100100101; end
            14'd4708 : begin out <= 64'b0010000111101000001001000110000000100111110101001010100010111010; end
            14'd4709 : begin out <= 64'b1010100101110010001010001101000110101001000110111010101011101001; end
            14'd4710 : begin out <= 64'b1010101110011100001001011100011100101010100100010010000010001101; end
            14'd4711 : begin out <= 64'b1010101000000010001001011110111100101010101110110010100110111100; end
            14'd4712 : begin out <= 64'b0010100000001000001010101111110110101001101010010010101011101000; end
            14'd4713 : begin out <= 64'b0010100000001110001000100111000000100010011001101001011011100011; end
            14'd4714 : begin out <= 64'b0010101110011010101010111010000010101001010010110010100011110101; end
            14'd4715 : begin out <= 64'b0010100110100010001010111110001110101000111110011010011111111100; end
            14'd4716 : begin out <= 64'b1001111100110111000111010010101000100001111101101010011100100100; end
            14'd4717 : begin out <= 64'b1010101011011001101001111010000010100000110111000010100100111011; end
            14'd4718 : begin out <= 64'b0010100110110000101010101101101110101000010000111010100110110011; end
            14'd4719 : begin out <= 64'b0010101110111001001000110000001100101001001010111010101110110110; end
            14'd4720 : begin out <= 64'b0001010011010001001010010010000010101001000000000010101111001000; end
            14'd4721 : begin out <= 64'b1001111110000011001001001010001010101010110100010010100100111111; end
            14'd4722 : begin out <= 64'b1010010110110101001010011010010110011011101000010010101101011010; end
            14'd4723 : begin out <= 64'b1010100111101010001010001010000010100111011001110010010010000111; end
            14'd4724 : begin out <= 64'b0010101011101000001001011101111100101001000001101010101011000011; end
            14'd4725 : begin out <= 64'b0010100100101001101010010110010110101001101001001000010000111010; end
            14'd4726 : begin out <= 64'b1010011100101100001010010001000010101010111000110010101000111001; end
            14'd4727 : begin out <= 64'b0010100010100101101010010010101100100101101101000010101101001110; end
            14'd4728 : begin out <= 64'b0010101100011101100110011011011000011110101110000010011110010101; end
            14'd4729 : begin out <= 64'b1010000000011111100110000001000000101010100001000010010101001000; end
            14'd4730 : begin out <= 64'b0010100001111001001010010001011110101011101111100010010011010100; end
            14'd4731 : begin out <= 64'b0010001100001000001001011110011010100010110110101010011010011001; end
            14'd4732 : begin out <= 64'b0010000110110000001010101010110010101011100010101010100111101001; end
            14'd4733 : begin out <= 64'b0010011000100010101010110101000010100011101000110010010110110010; end
            14'd4734 : begin out <= 64'b1010101111011111101010010011010110101001111011000010011111100100; end
            14'd4735 : begin out <= 64'b1010011111010100001010011100010000100010100010101010101110001011; end
            14'd4736 : begin out <= 64'b0010101011000110001010011110011000101000111110100001101000101101; end
            14'd4737 : begin out <= 64'b0010011010100000101001010000010010101001001011111010011011101000; end
            14'd4738 : begin out <= 64'b0010000001010011001010011001100010101010111101001010100010011011; end
            14'd4739 : begin out <= 64'b0010101000010100001010010111001110101001111010000010000001001101; end
            14'd4740 : begin out <= 64'b0010100010110000001010111001111010100100111011100010100111111001; end
            14'd4741 : begin out <= 64'b1010010011110001001000011110100100101100000101011010101101101010; end
            14'd4742 : begin out <= 64'b1010101000100001101010011011101000101000001110101010001111100110; end
            14'd4743 : begin out <= 64'b1010001001101101101001001000110110100010000010001010010101011000; end
            14'd4744 : begin out <= 64'b1010000011001101101000111100011010101000101000101010101000101001; end
            14'd4745 : begin out <= 64'b0010011111100110001010001011100100101010011111011010010000010001; end
            14'd4746 : begin out <= 64'b1010101110011001101010000100101110101001010111101010101000110011; end
            14'd4747 : begin out <= 64'b1010101110000110001000011101010110101011001100011010100100110010; end
            14'd4748 : begin out <= 64'b1010101100100001001000110111111110100111001101111010100100111010; end
            14'd4749 : begin out <= 64'b0010100010101100001000110011110110100100110010001010011110100111; end
            14'd4750 : begin out <= 64'b1010101111010000001010111000001010100111000111000010100001111001; end
            14'd4751 : begin out <= 64'b0001010110111111100111101100001000100101011110000010101111000110; end
            14'd4752 : begin out <= 64'b1001011000010111001001001000100110101011111011101010000000111110; end
            14'd4753 : begin out <= 64'b1010101011100111101010100001110000101000100000101010011100001101; end
            14'd4754 : begin out <= 64'b1010100010000111000111101010000100101001101010010010100011111100; end
            14'd4755 : begin out <= 64'b1010110001001010001001011110110100100100010111001010101100100100; end
            14'd4756 : begin out <= 64'b1010100000101111001000010101001110101001010011100010000001010011; end
            14'd4757 : begin out <= 64'b1010010110010110101010110101000010101001001001100010000101101110; end
            14'd4758 : begin out <= 64'b1010001011001011101010001101110000011101000110100010100011011100; end
            14'd4759 : begin out <= 64'b0010100010110011101000010111010000100101011010001010011101101011; end
            14'd4760 : begin out <= 64'b1010011100101010101001100110101000100000101001001001100000000011; end
            14'd4761 : begin out <= 64'b1010101110001011100010110110000100100110010101100010001011101010; end
            14'd4762 : begin out <= 64'b0001110101111100001010000101111000011111010100101010001000101100; end
            14'd4763 : begin out <= 64'b1010011100010101001010001011010000101011011000100010000101111000; end
            14'd4764 : begin out <= 64'b0010001011001001001000011101100000101011100101101010100101011100; end
            14'd4765 : begin out <= 64'b1010011001110010101010111100011000101011100101010010011011011100; end
            14'd4766 : begin out <= 64'b1010101110110000101001100100001010101001101010000010101011011110; end
            14'd4767 : begin out <= 64'b0010101111001000001000111000000100101000011101001010001101010001; end
            14'd4768 : begin out <= 64'b0010101011110011001010110001000000100101010101111001111000101010; end
            14'd4769 : begin out <= 64'b0010011101000110001010111001111010100011111100010010011101110001; end
            14'd4770 : begin out <= 64'b0010001110110101001010001001110010101010000000110001110110010111; end
            14'd4771 : begin out <= 64'b0010011100101100101001010010111010010010111101000010010100001111; end
            14'd4772 : begin out <= 64'b1001111010001100001001000000001000101011011100001001110001100011; end
            14'd4773 : begin out <= 64'b1010100101011100001010010101010000100110100011010010100101001100; end
            14'd4774 : begin out <= 64'b1010010010101111101001100100011010100100110010001010100100011110; end
            14'd4775 : begin out <= 64'b1010100111111001001010111110111110100011010000011010100001110000; end
            14'd4776 : begin out <= 64'b0001101111001000001010010000111010100111011101010010010001110100; end
            14'd4777 : begin out <= 64'b0010100001001001001010000100000110100011000000000010100101100100; end
            14'd4778 : begin out <= 64'b0010101101100100000111011011101000101001010101110001111001110011; end
            14'd4779 : begin out <= 64'b0001011011111000000111010011011000101000011110010001110011110001; end
            14'd4780 : begin out <= 64'b1010011011100000101010001010001000101000111011011000111100001010; end
            14'd4781 : begin out <= 64'b1010100011000110001010001101000010011011011101111010101000000010; end
            14'd4782 : begin out <= 64'b0010001010011001101001000010000010101000111110001010010111110010; end
            14'd4783 : begin out <= 64'b1010101001011101101010111011011110101001100011001001111000010100; end
            14'd4784 : begin out <= 64'b1001110001001011101001111010000110101010101001101010101101000100; end
            14'd4785 : begin out <= 64'b1010010011101111000110001000111110100100010100010010100100001011; end
            14'd4786 : begin out <= 64'b0010011001110010001000110011010010100001111111010001010001101001; end
            14'd4787 : begin out <= 64'b0010011100111100101010010101110000101011000011001010011110101010; end
            14'd4788 : begin out <= 64'b1010100010010000001010101101111110101000001010001001100101100011; end
            14'd4789 : begin out <= 64'b0010010111011011001010100101001000100101011111010010011101101110; end
            14'd4790 : begin out <= 64'b1010101010011100001010011001010100100011011011011010011000000111; end
            14'd4791 : begin out <= 64'b1010010110101110001010001011111010011001001110000010100000001101; end
            14'd4792 : begin out <= 64'b0010100110001001101010111010110010101011000100011010101000111001; end
            14'd4793 : begin out <= 64'b1010000001001000001010111110010100100110111000111010000000011000; end
            14'd4794 : begin out <= 64'b1010011111001100001000011100010110101011010111000010011101010011; end
            14'd4795 : begin out <= 64'b0010101110111010101010110110000100100011100100111010010111110110; end
            14'd4796 : begin out <= 64'b0010101100011001001001000111111110100100111110001010000010000011; end
            14'd4797 : begin out <= 64'b0010011101110000001010100001000000100100101100011010101110101110; end
            14'd4798 : begin out <= 64'b0010101001010110001010111011011000101001111101111010101111100000; end
            14'd4799 : begin out <= 64'b0010101001111110001010010100010110100000010101111010011010000111; end
            14'd4800 : begin out <= 64'b0010100000110010101001010011001010101000010011101010100101110100; end
            14'd4801 : begin out <= 64'b0010010110111011101010000100111000011111000111111010000100101101; end
            14'd4802 : begin out <= 64'b0010100010010101001001100111111100100011011010101010011010011111; end
            14'd4803 : begin out <= 64'b1010011001010100001010000100011000101011111011100001110000001100; end
            14'd4804 : begin out <= 64'b1010010101010011101010100101100010100101111100110010100000101111; end
            14'd4805 : begin out <= 64'b1010101111001011001001101101011100101011001010000010100001111100; end
            14'd4806 : begin out <= 64'b0010100111111100001000011101010010101000111110100010010110010110; end
            14'd4807 : begin out <= 64'b0010010000001010001010010010000000101000001100111001110000011001; end
            14'd4808 : begin out <= 64'b0010001111101110000111011111001110100110011000110001111010101011; end
            14'd4809 : begin out <= 64'b0010011011100101101000010011100000100100001101011010010000000011; end
            14'd4810 : begin out <= 64'b1010101111011001001001111111011110100110110101101010001100000010; end
            14'd4811 : begin out <= 64'b1010100001100100001010110010111100101010011110011010011101001101; end
            14'd4812 : begin out <= 64'b1010101110111001101001110111110010100111110011101001100011110000; end
            14'd4813 : begin out <= 64'b0010010010110100001001111110001000100111010111111010010111101000; end
            14'd4814 : begin out <= 64'b0010101110101000101001110001011010101001010100001010101011011010; end
            14'd4815 : begin out <= 64'b0010100100111011001001010001110000100100000100010010101101011110; end
            14'd4816 : begin out <= 64'b1010101111011010001000110100110000100111010100101010011110100111; end
            14'd4817 : begin out <= 64'b0010011000101111100110111000011110101010111000011010100100110100; end
            14'd4818 : begin out <= 64'b0010110001100000101010001000001100100011011101000010001101000011; end
            14'd4819 : begin out <= 64'b1010101010110110001001101110101100100100001000011010100000110000; end
            14'd4820 : begin out <= 64'b1010000101001110100110011111110010100010101100011010100011100101; end
            14'd4821 : begin out <= 64'b0010011001010111000110000001111000100100100011110010101100011100; end
            14'd4822 : begin out <= 64'b0010011101101010101001011100101010100110011001001010100111010101; end
            14'd4823 : begin out <= 64'b1010100011110100101001010001100100101000011100000010101010000110; end
            14'd4824 : begin out <= 64'b0010101100110001001001110010110100101010101010101010100011011110; end
            14'd4825 : begin out <= 64'b1010001010011000001010011011111000100110000001010010100001100000; end
            14'd4826 : begin out <= 64'b0010100000001001101001110001010010101011001010100010010001111100; end
            14'd4827 : begin out <= 64'b1010101011110001001001000110001110100110111010001010010110110001; end
            14'd4828 : begin out <= 64'b0010101010110010001010111000000010100011011001001010001100100010; end
            14'd4829 : begin out <= 64'b1000111100010111101010110111000000100100010110011010011000000101; end
            14'd4830 : begin out <= 64'b0010001111000011001010100101111110100101100011010010011110110011; end
            14'd4831 : begin out <= 64'b0010011010110100001010111011010000101010010001001010101100000110; end
            14'd4832 : begin out <= 64'b0010100100100101001010100000100000101001011000111001111111111111; end
            14'd4833 : begin out <= 64'b0010101010011101001001011001100010100111000011110010101011111100; end
            14'd4834 : begin out <= 64'b0010100110010111101010001011001110011100110011100010101001010011; end
            14'd4835 : begin out <= 64'b1010010000011010001000110001010010101010010110101010101001010110; end
            14'd4836 : begin out <= 64'b0010100110000011100111011110001000100100011101100010010110001010; end
            14'd4837 : begin out <= 64'b1010011011001000001001001010100010101010101101000010010100100100; end
            14'd4838 : begin out <= 64'b1010100001100011001001010001111110010100011110001010100110100010; end
            14'd4839 : begin out <= 64'b0010101001110000001001111100001010100101011000001010100011101111; end
            14'd4840 : begin out <= 64'b1010011000000110001001010001101100101001011011001010011011001101; end
            14'd4841 : begin out <= 64'b0010100111000110101010110001111100101000100000101010011101010111; end
            14'd4842 : begin out <= 64'b0010000111000001001010110101100110101000000001111010101001100011; end
            14'd4843 : begin out <= 64'b1010011000000101101001111111111010101011101101101010101100010101; end
            14'd4844 : begin out <= 64'b0000111110000110000111010001000100100001010000111010100101100011; end
            14'd4845 : begin out <= 64'b0010101111111110001001010010000110101011001100110010010100011001; end
            14'd4846 : begin out <= 64'b1010101111111100001000010111101010101000010001100010101001010010; end
            14'd4847 : begin out <= 64'b0010101101101101101010011101001010100101011011001010100001111101; end
            14'd4848 : begin out <= 64'b0010010101101111101010101010110010100101110010001010011100100010; end
            14'd4849 : begin out <= 64'b1010100101010111000110110000001100101011010000011010100000101010; end
            14'd4850 : begin out <= 64'b0010101100111110001010100100111110101001101101111010010011111110; end
            14'd4851 : begin out <= 64'b1010100110001110001001001101011010101001010001010010010010001100; end
            14'd4852 : begin out <= 64'b0010100100111110101001001001010110100101101001111010011100010101; end
            14'd4853 : begin out <= 64'b0010011011111000000111010011000010101011101101100010101110100110; end
            14'd4854 : begin out <= 64'b1010101010110110000111010000001100101001110001001010100111010001; end
            14'd4855 : begin out <= 64'b1010100001110000001010000001110100100111100010001010100101010101; end
            14'd4856 : begin out <= 64'b0010101100100110101010100001111010101011011001000010101110010011; end
            14'd4857 : begin out <= 64'b0010101101101100100101001101110000101000010011110010000111101101; end
            14'd4858 : begin out <= 64'b1010010010011100101010101111110100101000000001010001110010000001; end
            14'd4859 : begin out <= 64'b1010011100110110001010001001101100101011101100010010100111110001; end
            14'd4860 : begin out <= 64'b1010011010010001001010111101010010011111010011000010100000001011; end
            14'd4861 : begin out <= 64'b1010000001101001001001011010000010101010000111100010010110101111; end
            14'd4862 : begin out <= 64'b1010101100000110100011111010010010101010101101110010001010101000; end
            14'd4863 : begin out <= 64'b1010000111101011001010011001111100100001101001010010001101101111; end
            14'd4864 : begin out <= 64'b0010000011001111101000001111101000100001101000100010010111010111; end
            14'd4865 : begin out <= 64'b1010101011010110101001001010110110100101000101010010100100110100; end
            14'd4866 : begin out <= 64'b0010011000001011101010101000010010011101100101101010011110101110; end
            14'd4867 : begin out <= 64'b0010101000011011001001001110000000100110000111100001110100000001; end
            14'd4868 : begin out <= 64'b1010011111000000101010011010101110100100001101101010101001100110; end
            14'd4869 : begin out <= 64'b0010001001000110001010100100011100101000110100110001101111001101; end
            14'd4870 : begin out <= 64'b1010100111000010101010000110000000100110000110101001011100111011; end
            14'd4871 : begin out <= 64'b1010101000000100101010000000111010100101111100000001011000010111; end
            14'd4872 : begin out <= 64'b1010101001110101001010100010110110100101000001010010100110000011; end
            14'd4873 : begin out <= 64'b0010101010001011101010000101001100101010000001110010100110110110; end
            14'd4874 : begin out <= 64'b1010101110100111001010000110111010100101100101001010001010101010; end
            14'd4875 : begin out <= 64'b0010101000010001001000111110001000100110110010110010100001100010; end
            14'd4876 : begin out <= 64'b1010100010101111001010100110101110101001000000010010010110111111; end
            14'd4877 : begin out <= 64'b0001111100000000101001100011001010101000111111001010001011011010; end
            14'd4878 : begin out <= 64'b1010011100100111101000110000101110101001100000101010010110000110; end
            14'd4879 : begin out <= 64'b1001110010011100001000111001111000101001111111001010010110110011; end
            14'd4880 : begin out <= 64'b1010101111001101101001010101110010011010110000011010000101010010; end
            14'd4881 : begin out <= 64'b0010000100011100101010000101011100101010100110001010100100010000; end
            14'd4882 : begin out <= 64'b0010100001010110101010110011010010101000000010011010011011101111; end
            14'd4883 : begin out <= 64'b1010100101010100101010110000011110100111111110101010000111101101; end
            14'd4884 : begin out <= 64'b0010100010010001001000000101011000101001010010111010101010011110; end
            14'd4885 : begin out <= 64'b1010100000100111001000010111011000101001011010011001011011010110; end
            14'd4886 : begin out <= 64'b1010001110010011101010100110101010101010111101111010000001101110; end
            14'd4887 : begin out <= 64'b1001111001101001101000000000111010100011011010110010100011001011; end
            14'd4888 : begin out <= 64'b1001011110111111101010011100100100100100101011001010100100001000; end
            14'd4889 : begin out <= 64'b0010101110001000001000110100010000100101100110000010100100100111; end
            14'd4890 : begin out <= 64'b0010010011110101001001011101101110011100000101111010100111000100; end
            14'd4891 : begin out <= 64'b0010000000110001001001001110000010101000001001101010010011001101; end
            14'd4892 : begin out <= 64'b0010011101101001101010010001100100100100100101000010100010111001; end
            14'd4893 : begin out <= 64'b0010100101000101001010000011011000100111101110111010010100010011; end
            14'd4894 : begin out <= 64'b0010101110011101101010011010000110101001000000100010011111001000; end
            14'd4895 : begin out <= 64'b1010010111000011001000001111110000100101011100001001100111110100; end
            14'd4896 : begin out <= 64'b0010000110000010001001100101111010100110111110000010010011001011; end
            14'd4897 : begin out <= 64'b1010100001101100100110101001100110101001001111101010100011100110; end
            14'd4898 : begin out <= 64'b1010010100101100001011000000000100101000010001100010100101101111; end
            14'd4899 : begin out <= 64'b0010101011011001001010111010110110101010001110011010100110100110; end
            14'd4900 : begin out <= 64'b0010010001010011000110100001010000100101000000001010010011011000; end
            14'd4901 : begin out <= 64'b0010100111101100001000001011100110100110100010100010010000011101; end
            14'd4902 : begin out <= 64'b1010011101101000001010100100001000101010000011010010010111001010; end
            14'd4903 : begin out <= 64'b1010010101011110001010001000101110101011101000001010101010100010; end
            14'd4904 : begin out <= 64'b1001110111001111101001100111100110100110111000011010011011011110; end
            14'd4905 : begin out <= 64'b0010100111110100001010001010001110011011100100101010011100101010; end
            14'd4906 : begin out <= 64'b0001110111010110101010111010110100101011010000111010100001000000; end
            14'd4907 : begin out <= 64'b0010100000110001001010110010110010101011100010111010011111111110; end
            14'd4908 : begin out <= 64'b0010001001101100001001101001111110010101100111110010100111010110; end
            14'd4909 : begin out <= 64'b1010101101111011101010001101010010101011100001111010100001000111; end
            14'd4910 : begin out <= 64'b0010100000110001100110101100010110100100111000001010011111100111; end
            14'd4911 : begin out <= 64'b1001111010010001100110001101011110100111111100011010100100010110; end
            14'd4912 : begin out <= 64'b1010010110000000100100010101100110101010011011010010010001110011; end
            14'd4913 : begin out <= 64'b0001101000100110101010100111110000011001100111100010011101000000; end
            14'd4914 : begin out <= 64'b0010101110000001001000111111000000100100010110001010101011010011; end
            14'd4915 : begin out <= 64'b1010100011111011101010111101110110100110111011000010100001110001; end
            14'd4916 : begin out <= 64'b0010000001100101001010110001101010101010011110000010101101000011; end
            14'd4917 : begin out <= 64'b0010011010111110001001001001110110101000010101010010001000110100; end
            14'd4918 : begin out <= 64'b0010100001111111101000001101011000101011100000111010011101010000; end
            14'd4919 : begin out <= 64'b1001101000100010101010011011011110100011011101000010011011000010; end
            14'd4920 : begin out <= 64'b1010100011011001001010101000010000101000101110111010000011100110; end
            14'd4921 : begin out <= 64'b0010010000101001101000101110000110100111110110011010101001011111; end
            14'd4922 : begin out <= 64'b1010100100010111000101011010111000101011011101000010000010100111; end
            14'd4923 : begin out <= 64'b1010000101000000101010100101000110101010111011010010101110001110; end
            14'd4924 : begin out <= 64'b1010100001011100001010101001000110100111110011011010100001000001; end
            14'd4925 : begin out <= 64'b1010010110000001101010001101100010100110011010000010100110011110; end
            14'd4926 : begin out <= 64'b1010100110110001001010011000000100100111110000111010100011110110; end
            14'd4927 : begin out <= 64'b0010100010011001001010001000010010101011100001100010100110010111; end
            14'd4928 : begin out <= 64'b0010100100110011100110000100000010100110001100101010010000000110; end
            14'd4929 : begin out <= 64'b1010100011100111101010010111010000101001111000000010101110100101; end
            14'd4930 : begin out <= 64'b1010101010000110001001010110010010100010001110011010100110111101; end
            14'd4931 : begin out <= 64'b0010010001010011001001001101001100100101000101100010001010001101; end
            14'd4932 : begin out <= 64'b1010100110011100100110101111101000101010110111100010010000001001; end
            14'd4933 : begin out <= 64'b0010010011101101000111001100110100100010101110101010011011110101; end
            14'd4934 : begin out <= 64'b1010011111011101101010111001111100101000010000000010101101011011; end
            14'd4935 : begin out <= 64'b0010011010110111101010110111110110101010101001001010101001110101; end
            14'd4936 : begin out <= 64'b0001110111110011101010010001010100101100000011100010100110110000; end
            14'd4937 : begin out <= 64'b0010011010010101101001111010111010010110010111101010010101001111; end
            14'd4938 : begin out <= 64'b0010101111010101101010111110110000100100010000001010101010110101; end
            14'd4939 : begin out <= 64'b1010101110001101000110111110111110100111100111000010101011010001; end
            14'd4940 : begin out <= 64'b1010101101011001001010011010011010101001111101110010000101100110; end
            14'd4941 : begin out <= 64'b1010011110110001001001010100001000100110001010101001110011011011; end
            14'd4942 : begin out <= 64'b0010101110000101001010000110010100101000100000101010100010100010; end
            14'd4943 : begin out <= 64'b1010100111000011101001001011011010011011100011110010000101011100; end
            14'd4944 : begin out <= 64'b0010100010001110100111010101110000101011010100111010000010001011; end
            14'd4945 : begin out <= 64'b0010101001010100001010011011110000100110100111000010010000101111; end
            14'd4946 : begin out <= 64'b1001101111010000101010011101100010101011100110011001111010101101; end
            14'd4947 : begin out <= 64'b0010100110010101001001011101001110001100010101011010100011100000; end
            14'd4948 : begin out <= 64'b0010011000011001101001010010101010100101111100010010010100011011; end
            14'd4949 : begin out <= 64'b0010100111011001100100100111011100100000001000110010100010011000; end
            14'd4950 : begin out <= 64'b0010001001110111001010100110110010011101101010101010101010100010; end
            14'd4951 : begin out <= 64'b1010101100111001001010101010010110101010011010000010100100000001; end
            14'd4952 : begin out <= 64'b0001101101111001001010110000101010101011000101010010010001111110; end
            14'd4953 : begin out <= 64'b0010000001010011101010010110101100100011001101110010100000000100; end
            14'd4954 : begin out <= 64'b1010100010011000101010101001101000101010011000100010000110101011; end
            14'd4955 : begin out <= 64'b0010101011110100101010011001100000101011100111111010101001111000; end
            14'd4956 : begin out <= 64'b0010010100001010101010011010110100101010110001001001110000101010; end
            14'd4957 : begin out <= 64'b0010101011111110101010011000010100011101101001100001111110011000; end
            14'd4958 : begin out <= 64'b1010010100111101001010110011110010100101111101111010001101010000; end
            14'd4959 : begin out <= 64'b1010101000000001101001101011101110101001101111110010101010010010; end
            14'd4960 : begin out <= 64'b1010001111100111101010101001110110101011100110001010100100101010; end
            14'd4961 : begin out <= 64'b1010100110101000001010100010011100100000110010000010101111100000; end
            14'd4962 : begin out <= 64'b0010010101111111001010000000111010100111110111110010101001100011; end
            14'd4963 : begin out <= 64'b0010100001100000001010110101110100100100010111010001011010110011; end
            14'd4964 : begin out <= 64'b1001111101010010101010101011100010100000010100101010000101111101; end
            14'd4965 : begin out <= 64'b1010011000011010001010011010001000100010010011101010100100001110; end
            14'd4966 : begin out <= 64'b0010101101001001101010000110001010011000101101010001110011000101; end
            14'd4967 : begin out <= 64'b1010100111011011101001001001010000101011000101101010010011111011; end
            14'd4968 : begin out <= 64'b0010000001011000001010100000010000101000101111001010010010101100; end
            14'd4969 : begin out <= 64'b1010100000000100001001100101000010101000100111101010100011000000; end
            14'd4970 : begin out <= 64'b0010010010110001001000011110100000101000111010110010011010110110; end
            14'd4971 : begin out <= 64'b1010101010100110000110001111111010101000111101000010101001011000; end
            14'd4972 : begin out <= 64'b1010011001100111001000100100101110010011101100000010100110100010; end
            14'd4973 : begin out <= 64'b1010001101000000100101001101101110101000101000110010100010011110; end
            14'd4974 : begin out <= 64'b0010011000011100100110011111111010100100111011001010000001100101; end
            14'd4975 : begin out <= 64'b0001111110011011101001001100100100101010101000101010010011011110; end
            14'd4976 : begin out <= 64'b0010001000110011001010110000111010101010111111001010101111011111; end
            14'd4977 : begin out <= 64'b1010101001111001001010010000010100100111011100101010101000011010; end
            14'd4978 : begin out <= 64'b0001110111100111001000011100100000011011010100011010010010010111; end
            14'd4979 : begin out <= 64'b1010101000001111001010110100011110101010110011010010001111011101; end
            14'd4980 : begin out <= 64'b1001110000000001101001001011111110101000010000001010011111111011; end
            14'd4981 : begin out <= 64'b0010011100001110101010010000010110101000100011110010001111111011; end
            14'd4982 : begin out <= 64'b0010100100101010001000000100100110100111001000110010100101110101; end
            14'd4983 : begin out <= 64'b1010101110111011101010110000110100101011011111100010010010000110; end
            14'd4984 : begin out <= 64'b0010010100110011101010101101110000101010011010010010101011011100; end
            14'd4985 : begin out <= 64'b0010011010101000001010011101001100101011100111100001110000111110; end
            14'd4986 : begin out <= 64'b1010001011000000001010011111111010101010101010001010100111000100; end
            14'd4987 : begin out <= 64'b1010011101000000001001011100101010101001110101001010100110111001; end
            14'd4988 : begin out <= 64'b1010010000100011001010010111010000101010010101011010011101000111; end
            14'd4989 : begin out <= 64'b1010101011111000100111100101100010100101000000010010100100110010; end
            14'd4990 : begin out <= 64'b0010011010000010101010100111001110100000110000001010101100000110; end
            14'd4991 : begin out <= 64'b1010100111010110000110000111000100100100011001100010011111111001; end
            14'd4992 : begin out <= 64'b0010010110101100001001000100001000101001010110100010101001100111; end
            14'd4993 : begin out <= 64'b0010100110010100000101011010100010101010110111110010010100110010; end
            14'd4994 : begin out <= 64'b0010101001111000001000100111100100101000111110000010101010111110; end
            14'd4995 : begin out <= 64'b1010101000111011101010000100000100100000011001011010101001011001; end
            14'd4996 : begin out <= 64'b1001011011001101101001000011110010101011100010101010010001011100; end
            14'd4997 : begin out <= 64'b1010100111100111000100110101010100101001110111010010101010000010; end
            14'd4998 : begin out <= 64'b0010100001011001001010111111110010100101111110011010100001110110; end
            14'd4999 : begin out <= 64'b0010101110010010101001001100111100100100010001011010000111101001; end
            14'd5000 : begin out <= 64'b0010101001000101001010101010101000011100111100110010011101001011; end
            14'd5001 : begin out <= 64'b1010100011011111001011000000110010100011011101011010101100011110; end
            14'd5002 : begin out <= 64'b1010010001011010101001010000000010011111010100011010010100001011; end
            14'd5003 : begin out <= 64'b0010100110111010101001010111010010101011101001010001000000011111; end
            14'd5004 : begin out <= 64'b1010100101100010000111000001101010101000011001100010101100000000; end
            14'd5005 : begin out <= 64'b1010101001110110100111010101010000101011010110100010101011101011; end
            14'd5006 : begin out <= 64'b1001110111010111000111110011111010101000110000011001111000100111; end
            14'd5007 : begin out <= 64'b1010000110101001101001001011110010101011011000000010100101001000; end
            14'd5008 : begin out <= 64'b0010101000111100001001101000111110100111110100010010010101001010; end
            14'd5009 : begin out <= 64'b1010000001001111101010110110110100100011011111000010100111000001; end
            14'd5010 : begin out <= 64'b0001111010011001001001110100010110101001100111011010011000100010; end
            14'd5011 : begin out <= 64'b1010010111010101001010010100011010101000101101100010011101000011; end
            14'd5012 : begin out <= 64'b0010100110000001101010011010000110100011110110111010100111001000; end
            14'd5013 : begin out <= 64'b1010001111001111101011000011100000011010001110110010100010001001; end
            14'd5014 : begin out <= 64'b1010000000000100001010100110000110101000001011111010010111010000; end
            14'd5015 : begin out <= 64'b0010011111011010101010111010011100100101100101110010100111101100; end
            14'd5016 : begin out <= 64'b0010000010100001101010011111000100011100100001011010100101110010; end
            14'd5017 : begin out <= 64'b0010100011111011100100011100011100010010101100011010000010111001; end
            14'd5018 : begin out <= 64'b0000110001000000001010000111100110101011000100111010100001010010; end
            14'd5019 : begin out <= 64'b1010100101101010101010010011001110101000010101001010011011000110; end
            14'd5020 : begin out <= 64'b1001110111010111101010110011110010101010010111110010011011001111; end
            14'd5021 : begin out <= 64'b1001111010001010001010000001010110101010111010010010100110000000; end
            14'd5022 : begin out <= 64'b0010101001111100001010010111000110011110100011101001110111010011; end
            14'd5023 : begin out <= 64'b1001100010001111101000100000010000011000001110011010101000110010; end
            14'd5024 : begin out <= 64'b1010101100011101100111110100111100101001101110100010100010011010; end
            14'd5025 : begin out <= 64'b0001000100111011101010100101110100101000110101100010001110001010; end
            14'd5026 : begin out <= 64'b1010100110001000001010100101111110010110100111011010011101001110; end
            14'd5027 : begin out <= 64'b0010101101011001000111011111111010101010010111001001110001001011; end
            14'd5028 : begin out <= 64'b0010011111100111101010001100100010101001001011101010011010000111; end
            14'd5029 : begin out <= 64'b0010010111111011001011000001100100011110011011111010001111001000; end
            14'd5030 : begin out <= 64'b0010011000010001101010111001010000100111101101100010001110010111; end
            14'd5031 : begin out <= 64'b0001111011010011101001000011111000101001111000011010001100101010; end
            14'd5032 : begin out <= 64'b0001001100001111101010110001111110100010000101001010101010101111; end
            14'd5033 : begin out <= 64'b1010010110001010100111101111010010101011011111100010010111100111; end
            14'd5034 : begin out <= 64'b1010010001111111101010110101100000100101000011001010101111110111; end
            14'd5035 : begin out <= 64'b0010101001000100001010001101001010100000011000100010010001011110; end
            14'd5036 : begin out <= 64'b0010100001011111001001111111110010100101000011001010101010110001; end
            14'd5037 : begin out <= 64'b1010000111111001001010110110000110100111010011011010100011110110; end
            14'd5038 : begin out <= 64'b1010011000101111001010101110100110100100010111010001110101010000; end
            14'd5039 : begin out <= 64'b1010010000001111101001111000011110100100011001110001110110010010; end
            14'd5040 : begin out <= 64'b0010101101000000001001011110010100101001100000000010011001111000; end
            14'd5041 : begin out <= 64'b0010100011010100101010001000011000101010010000110010101101110101; end
            14'd5042 : begin out <= 64'b0010001110111111000111010001110110101011010010010010101010011100; end
            14'd5043 : begin out <= 64'b1010001111011101101010010100100010101000110101000010100001001000; end
            14'd5044 : begin out <= 64'b1010011100000000101000101011011100011001010001010001110001101011; end
            14'd5045 : begin out <= 64'b0001011000001001001001011100000010100111100100101001110010101111; end
            14'd5046 : begin out <= 64'b1010101001000001100111111111000000100110001111101010010111101100; end
            14'd5047 : begin out <= 64'b0010100010010100101010101000000010100100111110001010100011101000; end
            14'd5048 : begin out <= 64'b1010100000010101101001011001010110010111111000011010101001100010; end
            14'd5049 : begin out <= 64'b1010011011011010001010010010011000100001100001100010101110110100; end
            14'd5050 : begin out <= 64'b1010101110110110000110011011101000100000110000010010100110110100; end
            14'd5051 : begin out <= 64'b1010101010111010101010011110011000101011011010011010101011110000; end
            14'd5052 : begin out <= 64'b0010011110110110001001011110111000101011101001001001100100100101; end
            14'd5053 : begin out <= 64'b0010010001100110001010010000011000101000101001011001111110011001; end
            14'd5054 : begin out <= 64'b0010100001001000101010010101011100010001001101100010100011010111; end
            14'd5055 : begin out <= 64'b0010100110111101101010000010111100101000001100001010101011010001; end
            14'd5056 : begin out <= 64'b1010001010100010001001000011001100101010100111001010010100001000; end
            14'd5057 : begin out <= 64'b1010101101101000001000100011111000101001010000011010101001011000; end
            14'd5058 : begin out <= 64'b1001110100100101001010010011100110010000111010000010100111100111; end
            14'd5059 : begin out <= 64'b0010000010101010101010110011011010101000010111100001110000011111; end
            14'd5060 : begin out <= 64'b1010101010000010100101111000100010100100111111011010000110011011; end
            14'd5061 : begin out <= 64'b1010011110110110101001101001101100101000010101011010101111101110; end
            14'd5062 : begin out <= 64'b1001110001101010001010110001111110101000100100000010101001100111; end
            14'd5063 : begin out <= 64'b1010100101110100101010010111010000101001001001010010100100111000; end
            14'd5064 : begin out <= 64'b1010001100000110101010000100000110101010000000110010001110111110; end
            14'd5065 : begin out <= 64'b1001111110000001101010010100101110101001101110010010100111101011; end
            14'd5066 : begin out <= 64'b0010100111100011001010001100100000100110111111010010101001100100; end
            14'd5067 : begin out <= 64'b0010101110001110001001001100000010101001101100110010000011101010; end
            14'd5068 : begin out <= 64'b1010100110001100101010011110001110100001011110100010101101111000; end
            14'd5069 : begin out <= 64'b0010100001000011101010001010010000101011111000110010101000010100; end
            14'd5070 : begin out <= 64'b1010100100011010101000111110000100010000101000101010011011000001; end
            14'd5071 : begin out <= 64'b0010100010000101001000001010100010101000000100100010010011010101; end
            14'd5072 : begin out <= 64'b1010000010011110101010000000111000011110010110100001111001111011; end
            14'd5073 : begin out <= 64'b1010101001101011101001101010010110100001001110010010001011001000; end
            14'd5074 : begin out <= 64'b0010100010100000001011000101111010001011000000100010001101001110; end
            14'd5075 : begin out <= 64'b0010100001001110101000001000100100101001001010100010101000101001; end
            14'd5076 : begin out <= 64'b1010000110111111001010101000101100100101001001111010101110011001; end
            14'd5077 : begin out <= 64'b0010010101001110001010111010011010101000000100100010000101000010; end
            14'd5078 : begin out <= 64'b1010001111010100001000011011111010100001010000010010001001010011; end
            14'd5079 : begin out <= 64'b1010101011011000101000000101000110101001000110001010000101001001; end
            14'd5080 : begin out <= 64'b1010011011110001001001000101011110101010000011000010100011010111; end
            14'd5081 : begin out <= 64'b1010010001111100001001110101000010101010100010010010010101110110; end
            14'd5082 : begin out <= 64'b1010011110011101101010111001111010011000100110000001110110000001; end
            14'd5083 : begin out <= 64'b1010100100000011001010011011100100101000111010101010010011011001; end
            14'd5084 : begin out <= 64'b1010010011001011101000011010100010011011110110100010010110110111; end
            14'd5085 : begin out <= 64'b0010011101011101101000001110111010101011011110011010001011000110; end
            14'd5086 : begin out <= 64'b0010101010110111100110110101101000100111011010100010101011011111; end
            14'd5087 : begin out <= 64'b1010101100001101101001110011100110101010010100101001100111011101; end
            14'd5088 : begin out <= 64'b1010010001101011001000010010101000100110011110110010100101111010; end
            14'd5089 : begin out <= 64'b0010100111011100001010000111000000101001001001000010101001010101; end
            14'd5090 : begin out <= 64'b1010001111011101101010000001001100001101010101010010100100111111; end
            14'd5091 : begin out <= 64'b1010101011110100101010000011010110010110101101011010011010000110; end
            14'd5092 : begin out <= 64'b1010100000101001101001011010011000101010011000000010101011001110; end
            14'd5093 : begin out <= 64'b0010100111101000101000111000101000100101010101011010100100010100; end
            14'd5094 : begin out <= 64'b1010101110100110001000110000100010100101101011000010100010000101; end
            14'd5095 : begin out <= 64'b1010000001000001101010110011001110100101011001001001111111111010; end
            14'd5096 : begin out <= 64'b1010010000101011001010010011101000100110010000101010100111110000; end
            14'd5097 : begin out <= 64'b1010101000110001100111000001001100100111111011001010100110001100; end
            14'd5098 : begin out <= 64'b1010100010011100001000110010110110010101100001011001110010101010; end
            14'd5099 : begin out <= 64'b0010001001110111001001100010010100101011101000100010100110111100; end
            14'd5100 : begin out <= 64'b1010100001100011001001111011001100101001100111111010101100011000; end
            14'd5101 : begin out <= 64'b1000110111001011001000001000111100100110000010101010100000011011; end
            14'd5102 : begin out <= 64'b1000100110010101101010111111100010101000000001111010011100010100; end
            14'd5103 : begin out <= 64'b0010010010110110101010110010001100101000110001010010101100100100; end
            14'd5104 : begin out <= 64'b0010100110111011001010000101000010101000001101011010101011101010; end
            14'd5105 : begin out <= 64'b1001110001110011001010001010000110100001000010101010010000001101; end
            14'd5106 : begin out <= 64'b0010011101000101101010110000111010101000000110100010100001001111; end
            14'd5107 : begin out <= 64'b1001111001000011000110110110100100100110011100100010101010111111; end
            14'd5108 : begin out <= 64'b0010011000110111101010011001001100101010000000110010100000110110; end
            14'd5109 : begin out <= 64'b0010010110101111001010111111111010100100010111000010101011100001; end
            14'd5110 : begin out <= 64'b1010010101001011101011000110101000010000110110000010000110010000; end
            14'd5111 : begin out <= 64'b1010101101000001101010111101110100101010110011000001111100001000; end
            14'd5112 : begin out <= 64'b0010101001100010001010100000110100100111100010100010011011010101; end
            14'd5113 : begin out <= 64'b0010100110100110001010010000110010101000110000010010011011101000; end
            14'd5114 : begin out <= 64'b1010010100011101001000100111000100101000011110011010100000101110; end
            14'd5115 : begin out <= 64'b0010000110110110101010101101011000101001111100010010101101011000; end
            14'd5116 : begin out <= 64'b0010100010011111101010001000011000101001001101000010010001011000; end
            14'd5117 : begin out <= 64'b1010101000110100000101101010100100101010111011111010101111011010; end
            14'd5118 : begin out <= 64'b1010011111111010000111100000100010100010000101101010011001010011; end
            14'd5119 : begin out <= 64'b1010011111100000001011000011101100101010000000001010001101110000; end
            14'd5120 : begin out <= 64'b0010011110101110101001111110110110011110100101100010001110000000; end
            14'd5121 : begin out <= 64'b1010001111111000101010111101100110101000101110000001011111101100; end
            14'd5122 : begin out <= 64'b0001110101011100000110001100000000100001100111110010101010101010; end
            14'd5123 : begin out <= 64'b1010101011101111001000111101100000101001100011110010101111101000; end
            14'd5124 : begin out <= 64'b1010101000101010100011011101001110101010001011111010100110111100; end
            14'd5125 : begin out <= 64'b0010100010010000001010111011111100100101110010101010010011000010; end
            14'd5126 : begin out <= 64'b0010010010111010001010011100101010101010000100000010101010010001; end
            14'd5127 : begin out <= 64'b1010100011100101000110101001100000101000111000010010101111001100; end
            14'd5128 : begin out <= 64'b1010100010001100101001000110100010101011001010010010101100111111; end
            14'd5129 : begin out <= 64'b1010100100101001001010000000111000101001010101011010000110100110; end
            14'd5130 : begin out <= 64'b0010001111101011001001010011111000101010101011011010100010011101; end
            14'd5131 : begin out <= 64'b1010100100111101101001000111111000100010110100110010101100101100; end
            14'd5132 : begin out <= 64'b1010011110110110101000101011100110011101101101101010101000111100; end
            14'd5133 : begin out <= 64'b0010100101011011001010100100001100101011110010010010011001001111; end
            14'd5134 : begin out <= 64'b0010101111111111001001101111101110100101110101011010101100111011; end
            14'd5135 : begin out <= 64'b1010100100111111001010100001111100101001011010111010010101000000; end
            14'd5136 : begin out <= 64'b1010100111011111001010000110110000101001110010011010100010000000; end
            14'd5137 : begin out <= 64'b0010100110001101001010100101010110101001011111101010011110101110; end
            14'd5138 : begin out <= 64'b0010010111101110000111100111111100101011101100011010100101110000; end
            14'd5139 : begin out <= 64'b1010101001110110001010111000110100101010110011000010100101110011; end
            14'd5140 : begin out <= 64'b1010101001100001001010101100011110001100010111011010010100000011; end
            14'd5141 : begin out <= 64'b1010100000001101101001010000000000100101010100010010101010000011; end
            14'd5142 : begin out <= 64'b0010101000000100101010011011100110011110100001110010101110100110; end
            14'd5143 : begin out <= 64'b1010100001000111001000111100111000101001100010101010100110011111; end
            14'd5144 : begin out <= 64'b1010101110000011001000001010001000100001000000001010100100000000; end
            14'd5145 : begin out <= 64'b0010001001110101101010011001011100101001111011110010001100000010; end
            14'd5146 : begin out <= 64'b0010101101010110101010011100101000101000101000110010100011110001; end
            14'd5147 : begin out <= 64'b0000010101011011101010010100001110101001011010011010001001110101; end
            14'd5148 : begin out <= 64'b0010101111000011101010101100110010101010010000011010010010110100; end
            14'd5149 : begin out <= 64'b1010010110111011001010100100110010101010011001010010000101010000; end
            14'd5150 : begin out <= 64'b0010011101111100000011101000111000100001010011101010100110110110; end
            14'd5151 : begin out <= 64'b0001110100001011101010100001110010101001001111110010101000100001; end
            14'd5152 : begin out <= 64'b1001111011001100101010100001001100100101110011111010101000101111; end
            14'd5153 : begin out <= 64'b1010010000000011001010101011011010101000111011010010011011110010; end
            14'd5154 : begin out <= 64'b0010101100100011101001001110011100100010001100011000111011101101; end
            14'd5155 : begin out <= 64'b0010011010011111001001101001010000101100001010010001110101100010; end
            14'd5156 : begin out <= 64'b0010100001001000001010110010100110101010000100100010101010110000; end
            14'd5157 : begin out <= 64'b1010101101101100001010010100001000100110010011011001100111000101; end
            14'd5158 : begin out <= 64'b0010001101101101101010011000101000101011100100011010101001111011; end
            14'd5159 : begin out <= 64'b1010011111010101101000111010110010101001000100111010010100100011; end
            14'd5160 : begin out <= 64'b0010010111100001101000100011010010101011011100000010010010111100; end
            14'd5161 : begin out <= 64'b1001101001001111101000111000001000011001010111110010011011000001; end
            14'd5162 : begin out <= 64'b1010000100010100000111011000110010101001000001011001110100101111; end
            14'd5163 : begin out <= 64'b0010100111100100101001011100010100101010000100110010100011101111; end
            14'd5164 : begin out <= 64'b1010100010010101100101011000001010100000101100011010100010100011; end
            14'd5165 : begin out <= 64'b0010101110011011001010100000001000100100010100110001110000100101; end
            14'd5166 : begin out <= 64'b0010011110000110001010111000001110101000100110011010100010011011; end
            14'd5167 : begin out <= 64'b0010101110110101101010110100110010100110001010001010100110011001; end
            14'd5168 : begin out <= 64'b1010100101111110001001000110011110101000110010010010011001111001; end
            14'd5169 : begin out <= 64'b0010100110110101001001110101010100101001000011001010000101001001; end
            14'd5170 : begin out <= 64'b1010101110000001101010100100100010101000011110111010100011111001; end
            14'd5171 : begin out <= 64'b0010001000011011001010001111000010101010011101001010001000110100; end
            14'd5172 : begin out <= 64'b1001110100010010101001000111010100100001110101111010001001011101; end
            14'd5173 : begin out <= 64'b1010010111100011101000110000011110011111110010100010010010001001; end
            14'd5174 : begin out <= 64'b0010011011000100101010000000111100101000001001011010101000010011; end
            14'd5175 : begin out <= 64'b0010011111000001101010011110001100100011111101010010100111100111; end
            14'd5176 : begin out <= 64'b1010010110101110101010011111010000101001001111111010100101001001; end
            14'd5177 : begin out <= 64'b0001100010100110000101111011011110100111001010001010100111100000; end
            14'd5178 : begin out <= 64'b0010011111001011001010010110010000100111110000111001101000110000; end
            14'd5179 : begin out <= 64'b0010011011101101000111000010111110101011000110010010001011001111; end
            14'd5180 : begin out <= 64'b0010011001110100001010011110001010100100111101101001001111010011; end
            14'd5181 : begin out <= 64'b0001110101100011001001001000110110101011110100100010100111101110; end
            14'd5182 : begin out <= 64'b1010000000011111101010110100100100100110101110010010101011110011; end
            14'd5183 : begin out <= 64'b1010100001010110001010111111011100101001010100010010101000100011; end
            14'd5184 : begin out <= 64'b0010100001101111101010100100100110101001100010001010011001010011; end
            14'd5185 : begin out <= 64'b0010101000101111101010100100111110101011101001110010011111011111; end
            14'd5186 : begin out <= 64'b0010011001001101101010110110111110001100011101011010011100101111; end
            14'd5187 : begin out <= 64'b0010100001101101101010100000101000101001101110011001011101001000; end
            14'd5188 : begin out <= 64'b1000101111000010000110000101001100101001101101111010100011100101; end
            14'd5189 : begin out <= 64'b1010101100110011001010011011100100101000000111111010100110100000; end
            14'd5190 : begin out <= 64'b1000111001101100101000111100010110100111100011001010100011111101; end
            14'd5191 : begin out <= 64'b1010001101110110001010000110110110100101101001001010100001110010; end
            14'd5192 : begin out <= 64'b1010100100100010001001001111001000011100011011101010101110101100; end
            14'd5193 : begin out <= 64'b1010101110001110101010010011110000100111000011110010001111110011; end
            14'd5194 : begin out <= 64'b0010100010001001001010011000101000101010101000111010010110110101; end
            14'd5195 : begin out <= 64'b1010100100101011001010101101011010010111110101000010100110100111; end
            14'd5196 : begin out <= 64'b0010101110101101101001101001000000101001110111001010100100000010; end
            14'd5197 : begin out <= 64'b0010001110010110101010101011001100101011100101111010101100100111; end
            14'd5198 : begin out <= 64'b0010010000110100101010011010101100011110010001001010001111011110; end
            14'd5199 : begin out <= 64'b0010101110001010101010010011111110101011101010100010100001101111; end
            14'd5200 : begin out <= 64'b1010001101000001001001000011100100101011011000011010100000111000; end
            14'd5201 : begin out <= 64'b1010100001001111101010011011011000101001000101010010100001011111; end
            14'd5202 : begin out <= 64'b1010101110001101001001011000001100101000000010100010011010010000; end
            14'd5203 : begin out <= 64'b0010100100011001001010000010001100100100001100111000100010010101; end
            14'd5204 : begin out <= 64'b0010100100101010101000100010000110100000111001101010101011111111; end
            14'd5205 : begin out <= 64'b1010100101101001001000011011111110101001111000101010100011111111; end
            14'd5206 : begin out <= 64'b1010100000101110001010110110001000101001100100011010010010000101; end
            14'd5207 : begin out <= 64'b0001100000000110001010111001010000101010101111110010100001110100; end
            14'd5208 : begin out <= 64'b1010010101100100101010000100100100011000111000110010100111110101; end
            14'd5209 : begin out <= 64'b0010011100111001000111001111110010100101010000000010101011000001; end
            14'd5210 : begin out <= 64'b1010100010011000101001011011110010100010001110000010101100001101; end
            14'd5211 : begin out <= 64'b1010000011001000001010011110100100011111011000111010101100000001; end
            14'd5212 : begin out <= 64'b0010000011111001001010101111000010100001010001011010001000111100; end
            14'd5213 : begin out <= 64'b1010000010111010001010101101000110100110111001111001010010001111; end
            14'd5214 : begin out <= 64'b1010000100001100001010101000001010101010000110000010101100010011; end
            14'd5215 : begin out <= 64'b0010100110110100101001001111001010100111111000011010010010011110; end
            14'd5216 : begin out <= 64'b1010011001001010001010010101101010100000111111010010011001000111; end
            14'd5217 : begin out <= 64'b1010100100001100001000110111010000100101010010101010010111100010; end
            14'd5218 : begin out <= 64'b0010100001100001001001010110111010100101011000010001110101110001; end
            14'd5219 : begin out <= 64'b1010000101110110001010011101100100011111110100111010010100000001; end
            14'd5220 : begin out <= 64'b1010101110011110101000100011111000011111011101010010010000000000; end
            14'd5221 : begin out <= 64'b1010101100011111001010101000000010101011001000011010100000001101; end
            14'd5222 : begin out <= 64'b0010000010100010101001001101111000100000000011001010001001100000; end
            14'd5223 : begin out <= 64'b0010101110100001101000011010111000101010101110110010010010011100; end
            14'd5224 : begin out <= 64'b1010010000110111101010110010101110100010010001111010010100100111; end
            14'd5225 : begin out <= 64'b0010011101111111001010000001010110101001110110010010100011101000; end
            14'd5226 : begin out <= 64'b1010101011000110001010110101001100100101110001101010011000011100; end
            14'd5227 : begin out <= 64'b1010100000101101001010011010001010101000111010001010101001111011; end
            14'd5228 : begin out <= 64'b1010101101101010101010101011100000101010011001000010010010100000; end
            14'd5229 : begin out <= 64'b1010011101101010001001000010110000101001110101101010011100110001; end
            14'd5230 : begin out <= 64'b0010001010100001100111110011110100100110100001011010101011101001; end
            14'd5231 : begin out <= 64'b0010101111111100100001100010000110101011110001010010100111010001; end
            14'd5232 : begin out <= 64'b1010010101000111101001110100000100101011101011100010100111100111; end
            14'd5233 : begin out <= 64'b1010010001001001101001110111010110011101011110000010100111110100; end
            14'd5234 : begin out <= 64'b1010010000110011101000011100000000101000101001010010101000111011; end
            14'd5235 : begin out <= 64'b1010100110101111001010111011011100101001110000101010100101100111; end
            14'd5236 : begin out <= 64'b0010001011111011101000100111010100101000101011111010100001011001; end
            14'd5237 : begin out <= 64'b1010100000001101101001110100010110100100010010111010101100110010; end
            14'd5238 : begin out <= 64'b0010011000100010101010001100100010101001001110001010000000101011; end
            14'd5239 : begin out <= 64'b1010100000100100001010101011101100101010110000011001011010000011; end
            14'd5240 : begin out <= 64'b1010101000100101001010011110100010100101100101011010101001010100; end
            14'd5241 : begin out <= 64'b0010101101011100001000100001101000101000110010011010011001011110; end
            14'd5242 : begin out <= 64'b1010100001111011101010001111101000100111010001111010100111111100; end
            14'd5243 : begin out <= 64'b1010011111101011100110010000101110100110111100011010101000010010; end
            14'd5244 : begin out <= 64'b0010100110100101001010010100100110101010100100110010100101100111; end
            14'd5245 : begin out <= 64'b0010101101011010101010010011010110101011110001111010100011111011; end
            14'd5246 : begin out <= 64'b0010100000000010001001010011110010011100000001010010011001010010; end
            14'd5247 : begin out <= 64'b1010011010101010100111000000110000100110000100000010101100011101; end
            14'd5248 : begin out <= 64'b0010100100011000001010001010000000101001110010111010010011101111; end
            14'd5249 : begin out <= 64'b0010000110110001001010111010111100101011101110001010001110010001; end
            14'd5250 : begin out <= 64'b0010000101001001001010001000001110101001100011100001110010011110; end
            14'd5251 : begin out <= 64'b0010110000011000101001011100010110100110101000001010100101000011; end
            14'd5252 : begin out <= 64'b1010101110001000101001110100110100101010010000110010110000000011; end
            14'd5253 : begin out <= 64'b1010101110011011001001101110000010011001001110111010101011111100; end
            14'd5254 : begin out <= 64'b0010100100101000000101000111000100101100010110001010100000111110; end
            14'd5255 : begin out <= 64'b0001001110011000001010001110110110100110011100001010100000101111; end
            14'd5256 : begin out <= 64'b0010011111011100001001110100110110100111000101001010011111011001; end
            14'd5257 : begin out <= 64'b1010101010011100001001111111111110100111101100001010100110110001; end
            14'd5258 : begin out <= 64'b0010101000011001101001011110010110011110101100111010011001001010; end
            14'd5259 : begin out <= 64'b1010101011110011101010011011100100100110111011100010001011110101; end
            14'd5260 : begin out <= 64'b0010101101011000101010110000010110101001001100110001100000111010; end
            14'd5261 : begin out <= 64'b0010100110110011001010010011110100101000100111101010011111100111; end
            14'd5262 : begin out <= 64'b0001110110000010101001000000011100101010010111111010100111100110; end
            14'd5263 : begin out <= 64'b1010010101010010101010001010111000101010110110010010101100010011; end
            14'd5264 : begin out <= 64'b0001010110010101001010010001010000100101111001100010011010100110; end
            14'd5265 : begin out <= 64'b1010010001110011001010100110111000101000010101101010000111010011; end
            14'd5266 : begin out <= 64'b1010010000101101000111010101110010100110100001111010101111111100; end
            14'd5267 : begin out <= 64'b0010010100011000101010000101001000100011010101111010100001101111; end
            14'd5268 : begin out <= 64'b1010100101111110001010011111010100101011100010001010011110110110; end
            14'd5269 : begin out <= 64'b0010011000111100001010010111110010100010000101100010000000110100; end
            14'd5270 : begin out <= 64'b0010000001001010101010100000010100101001111011111010101001000001; end
            14'd5271 : begin out <= 64'b1010100010001111001010100100010110100111100000101001001001110101; end
            14'd5272 : begin out <= 64'b0010011001001100101010000101101010101011110111011001111100001010; end
            14'd5273 : begin out <= 64'b0010000011000101001000010010010110101000000100100010100011101001; end
            14'd5274 : begin out <= 64'b1010011010100100001001011101000110101001111100100001101011100111; end
            14'd5275 : begin out <= 64'b0010101111010000001010001101101100100101001110000010011001011000; end
            14'd5276 : begin out <= 64'b1010000011101111101010111100110000100100001011000010101011000001; end
            14'd5277 : begin out <= 64'b0010100011110101001010001101011000011101011111100010101001111010; end
            14'd5278 : begin out <= 64'b1010100010000110101001000101110000101000101010001010101111011000; end
            14'd5279 : begin out <= 64'b1010001111100011001001001111110000101001100101010010101000011010; end
            14'd5280 : begin out <= 64'b1010010110101101101010010101110110011011111101111010000111011101; end
            14'd5281 : begin out <= 64'b0010101010000001000111101111011110100101000101001010011001010101; end
            14'd5282 : begin out <= 64'b1010101010111011001000010010000010101011001000111010100110000000; end
            14'd5283 : begin out <= 64'b1001100010100100101010001011001100100111111111000010001101011110; end
            14'd5284 : begin out <= 64'b1010011011000001100111111010110000100011110011100010101010111101; end
            14'd5285 : begin out <= 64'b0010100101111100101010010110100110010101111100011010101000000111; end
            14'd5286 : begin out <= 64'b1010100000101100001010111000001100101000101010011010100100111010; end
            14'd5287 : begin out <= 64'b1010100000001100001001001011000000101010110110000010011111010001; end
            14'd5288 : begin out <= 64'b1010110000001101101010100000111000101001001011011010001111001111; end
            14'd5289 : begin out <= 64'b1010011101001101001001011001011100101000101110001010010111111111; end
            14'd5290 : begin out <= 64'b1010101000001011001000000111101110011110111110010010101101000001; end
            14'd5291 : begin out <= 64'b1010100010000101001010100110110100011101011001100010010011000001; end
            14'd5292 : begin out <= 64'b0010101010000110001001000101011100101011011100110010100101001101; end
            14'd5293 : begin out <= 64'b0010100100001110001001011000100100101011000110101010100101101001; end
            14'd5294 : begin out <= 64'b0010101100101001001001101111000010011100111101011010100101101100; end
            14'd5295 : begin out <= 64'b1010000010001011001001000110000010101011011000010010101000111111; end
            14'd5296 : begin out <= 64'b0010000000001110100110000011000010011110000000101010011000110111; end
            14'd5297 : begin out <= 64'b1010100110000001001010100011011000100111100010010010010010010001; end
            14'd5298 : begin out <= 64'b1010100001000001101010100000101000101010010111101000010101111000; end
            14'd5299 : begin out <= 64'b1010110000000011001010011000011100100111011111000010011100001111; end
            14'd5300 : begin out <= 64'b1010101001000010001001100101001000101000010101101010100101100011; end
            14'd5301 : begin out <= 64'b1001100010000111101010000111111000011100111111001010101010100100; end
            14'd5302 : begin out <= 64'b0010101101001010101000111100011110100110001010111010100001101000; end
            14'd5303 : begin out <= 64'b1010011100110110101010000101010100101001100000011001111011001101; end
            14'd5304 : begin out <= 64'b0010001100110101001001100001011100011101000001110010100101100111; end
            14'd5305 : begin out <= 64'b1010100100101010101010010010001010100111011010011010100000100111; end
            14'd5306 : begin out <= 64'b1010011001110010101000011011010000011111111000010010000011001111; end
            14'd5307 : begin out <= 64'b0001101011010000001001110111010010011000110010001010100111010110; end
            14'd5308 : begin out <= 64'b1001101001111001100001111111100010100101110000100001001110001011; end
            14'd5309 : begin out <= 64'b1010010011000110100110100010011000100100100001111010100100010101; end
            14'd5310 : begin out <= 64'b0010101101001100101010100000100010100011011111011010100101000010; end
            14'd5311 : begin out <= 64'b1010101001100011101010011101010100101000101110001010011100111001; end
            14'd5312 : begin out <= 64'b0010100001001010001001111010011100100001111010011010101010000001; end
            14'd5313 : begin out <= 64'b0010101101011101001010101101011010101001110010111010001111111100; end
            14'd5314 : begin out <= 64'b0010101101010011001010111111000000101011010101000010100000101100; end
            14'd5315 : begin out <= 64'b1001110001110011001001000101100000100101100110111010101000000100; end
            14'd5316 : begin out <= 64'b1001110011011011101001011011110000101001100011100001110000111100; end
            14'd5317 : begin out <= 64'b1010010100010001001001001000000100100001100110011010101101100011; end
            14'd5318 : begin out <= 64'b0010011011101000000101100101100000011001011101001010101010000110; end
            14'd5319 : begin out <= 64'b0010011001111010101010111111010100101001101011011010100111001011; end
            14'd5320 : begin out <= 64'b1010101011010001101001111011111100101000101010010010101110011010; end
            14'd5321 : begin out <= 64'b0010101100110010001010101110011010101000110101001010001110100100; end
            14'd5322 : begin out <= 64'b1010100011110110001010100010010100011111010101100010010000010000; end
            14'd5323 : begin out <= 64'b1001110101001101101000101110000000011001101100101010000111011110; end
            14'd5324 : begin out <= 64'b1010101010101100001010000011101000101010110010010001110011101110; end
            14'd5325 : begin out <= 64'b1010100000010101001010100010011100101001101011100010101110100100; end
            14'd5326 : begin out <= 64'b0010010010100000101000111111001100011101010111000010101001000110; end
            14'd5327 : begin out <= 64'b0010100010011001101000000111001110101010111010101010101000001101; end
            14'd5328 : begin out <= 64'b1001111100000011101010100011001110101010011111110001101011010111; end
            14'd5329 : begin out <= 64'b1010101010010110101010001001101110011001000101011001111100000110; end
            14'd5330 : begin out <= 64'b0010011111011001001010001001010010011101001010111010010001111100; end
            14'd5331 : begin out <= 64'b1010011101101100100101000110101100100011010101010010100100000101; end
            14'd5332 : begin out <= 64'b0010101100000111101001010110010010101011010111010010011100101000; end
            14'd5333 : begin out <= 64'b0001101101101101000101101110001000101001110111100010011111111001; end
            14'd5334 : begin out <= 64'b0010101010111100001010001001110110101000101001111010001000000110; end
            14'd5335 : begin out <= 64'b0010011000101101000101000011101010100010001110110001100010101101; end
            14'd5336 : begin out <= 64'b1010011100101000001001101111010110100100001101110010011010100100; end
            14'd5337 : begin out <= 64'b1001101100000110001000111010100000101001010100001010101001111000; end
            14'd5338 : begin out <= 64'b0010010110110010001001001100101100101011010011110010101011010001; end
            14'd5339 : begin out <= 64'b0010011110001110101010000110100100100111111000111001011111000011; end
            14'd5340 : begin out <= 64'b1001110011000101001010000010111000100101100111110010011011111011; end
            14'd5341 : begin out <= 64'b0010100101011010101010010010110000011101001011010010010011101110; end
            14'd5342 : begin out <= 64'b1010100001000110001010101111001000101001111111111010010011011100; end
            14'd5343 : begin out <= 64'b1010001000010100101000011010001000101011011101100010101001010110; end
            14'd5344 : begin out <= 64'b1010101001101100001010000110001000011110101000100010010100010000; end
            14'd5345 : begin out <= 64'b1010011110100101001001101100110100011010010110111010010101000001; end
            14'd5346 : begin out <= 64'b1010100011010010000111010100111100101001011001110010010010001101; end
            14'd5347 : begin out <= 64'b1001111001011010101010010001110100100110010100111010101000000111; end
            14'd5348 : begin out <= 64'b1010010000100111001000111001001110101000100000100010000100110011; end
            14'd5349 : begin out <= 64'b0010101001011011001010100110101110100111101010000010001101000010; end
            14'd5350 : begin out <= 64'b1010011001101111101001110001111010100000101100101010101001100101; end
            14'd5351 : begin out <= 64'b0010100000111000101010111110000010101011110110100010101000111111; end
            14'd5352 : begin out <= 64'b1010100001111000101010101101001010101011010110101010010000011101; end
            14'd5353 : begin out <= 64'b0010010011011111101001111100011010100100010101011010100100010001; end
            14'd5354 : begin out <= 64'b0010010101101110001010011101010100101010110010100010101001010001; end
            14'd5355 : begin out <= 64'b0010011001010011101001000101111000101010101101001010110000001101; end
            14'd5356 : begin out <= 64'b1010011111110110001001011010000110101011011101111010010010001000; end
            14'd5357 : begin out <= 64'b0001111111000011001000001101110010101011001110001010010100011110; end
            14'd5358 : begin out <= 64'b0010010101010100100111110101000000100001111001111010100101111110; end
            14'd5359 : begin out <= 64'b1010101010100001101010001101001110101011001000011001110000011010; end
            14'd5360 : begin out <= 64'b0010101010111111101000000000011100101011001100011010001000010010; end
            14'd5361 : begin out <= 64'b0010100111001111001000010010001100101000000110001010100100011110; end
            14'd5362 : begin out <= 64'b1010000100000100101001000101111010101000110100000010100101100010; end
            14'd5363 : begin out <= 64'b0001111100111101001001010011111000100110111101101010011110000110; end
            14'd5364 : begin out <= 64'b0001100010100000001001001011011110100100011111010010010110011110; end
            14'd5365 : begin out <= 64'b0010000110001100101010010010100100101010010100010010101000111000; end
            14'd5366 : begin out <= 64'b1010010100011110101001011101100000101000000010101010101000100101; end
            14'd5367 : begin out <= 64'b0001111000110000101010111100011100101011101100010010101000110000; end
            14'd5368 : begin out <= 64'b0010010000000000001010010001101110101011111100010010101100000101; end
            14'd5369 : begin out <= 64'b0010100100101010101010101111011010101001100001011010001010111010; end
            14'd5370 : begin out <= 64'b0001111110001100001001011001100000100111101011010010001100001000; end
            14'd5371 : begin out <= 64'b0010011001100011101001000101101010011100100011010010001001101110; end
            14'd5372 : begin out <= 64'b0010011001000001001010100100001010101000011001010001101111000000; end
            14'd5373 : begin out <= 64'b1010100010010110101000101011111100101011011010001010101111111010; end
            14'd5374 : begin out <= 64'b1010000100111000001010011010011110011110100000101001100101111010; end
            14'd5375 : begin out <= 64'b0010100010010011101010101110000000101100010011111010100100100010; end
            14'd5376 : begin out <= 64'b1010000111001011001010010000001100100001101010111010100010111110; end
            14'd5377 : begin out <= 64'b0010101010000011001010111011010010101001001000101010101010101111; end
            14'd5378 : begin out <= 64'b1010101111110110101000011100000110000111000110110010101101001101; end
            14'd5379 : begin out <= 64'b1010100111000110001010010100011000101011011110110010101011001100; end
            14'd5380 : begin out <= 64'b0010100111010101101010001100101110101000111010111001111111011110; end
            14'd5381 : begin out <= 64'b1010100001100010101011000001100110011110010110010010101011001000; end
            14'd5382 : begin out <= 64'b0010101001111001101010101010111010100100100101111001101100111100; end
            14'd5383 : begin out <= 64'b1010101000001011001001010001010110010001110110000010101111010010; end
            14'd5384 : begin out <= 64'b0010100101111010101010000010000000100110010010100001111010000100; end
            14'd5385 : begin out <= 64'b1010100100110001101001011111101110100000000100100010011010000010; end
            14'd5386 : begin out <= 64'b1010101100001101101000000111000000011100010000110001110000100001; end
            14'd5387 : begin out <= 64'b1001111000011001101001110010111110101000101010101010101110011001; end
            14'd5388 : begin out <= 64'b0010100111010010101000010110111010101000101100001010001100101000; end
            14'd5389 : begin out <= 64'b1010100001111111001001011010010000011000010100100010100110101000; end
            14'd5390 : begin out <= 64'b0010010110100011001001101001010110011110010011100010000010010010; end
            14'd5391 : begin out <= 64'b0010101000000000001010111000010100100111111101001010011101010101; end
            14'd5392 : begin out <= 64'b0010101110111001100111110010101000011110100010011010010010001011; end
            14'd5393 : begin out <= 64'b0010001001010010001010011010110010100100111111111010100000000111; end
            14'd5394 : begin out <= 64'b1010100010011010101010101000110110101001101100010010100010010101; end
            14'd5395 : begin out <= 64'b0010000111010110101010001111000010100101111010110010010111011011; end
            14'd5396 : begin out <= 64'b1010010000011111101001110111111100101011100110100010001010101110; end
            14'd5397 : begin out <= 64'b1010011111100111101010010001001110100101100000010010101010001111; end
            14'd5398 : begin out <= 64'b0010101101101010101001011101011000100010100111001010101111011010; end
            14'd5399 : begin out <= 64'b1010010011000010101010100101110000100100001101010010010111110100; end
            14'd5400 : begin out <= 64'b0010101100100000100110101000001000100110111001010010000001011010; end
            14'd5401 : begin out <= 64'b0010010101011110101001110101000000100000111111001010100001001000; end
            14'd5402 : begin out <= 64'b0010110000000100001001000000001100101011001011110010011000011110; end
            14'd5403 : begin out <= 64'b0010100010110101000111001001001110101011101000101010101000001101; end
            14'd5404 : begin out <= 64'b0010010000101101001010010111100000101000011010000010011111111010; end
            14'd5405 : begin out <= 64'b0001100110001011001001101111010000100110111110111010101001101100; end
            14'd5406 : begin out <= 64'b1010011111100000001010000100010010011001010110100010000101010011; end
            14'd5407 : begin out <= 64'b0010101011101010101001100000110110101001000010000010100101010000; end
            14'd5408 : begin out <= 64'b1010010001010010001010001000110100100110011011010010100100101101; end
            14'd5409 : begin out <= 64'b0010100001111010101010101001111110100011100000010010100100011001; end
            14'd5410 : begin out <= 64'b0001000110100010100100110001001000100101101100010010000001000101; end
            14'd5411 : begin out <= 64'b1010100000000110001001101100110110011100000010010010011101011110; end
            14'd5412 : begin out <= 64'b0010101100101001001010111011001000010001111011010010100001110011; end
            14'd5413 : begin out <= 64'b0010101100011011001001100101000110100100000011110010011101110001; end
            14'd5414 : begin out <= 64'b1010101011011001101001101011001110101010011110000010100010001101; end
            14'd5415 : begin out <= 64'b1000110011110111100111000111010100101011011111100010010001100101; end
            14'd5416 : begin out <= 64'b0010101010111011001010110001011110100010100010111010010111010001; end
            14'd5417 : begin out <= 64'b1010010111001110000111110110000110100110100100111010101100000010; end
            14'd5418 : begin out <= 64'b0010100110111101001000000001110110101000101010100010100011011101; end
            14'd5419 : begin out <= 64'b1010101101101111101001101001101010011100100011111001111011011110; end
            14'd5420 : begin out <= 64'b0010010011100110101001100001111100101000111100101010000101011010; end
            14'd5421 : begin out <= 64'b0010100000010100101010111000100000101000001110001010101110110010; end
            14'd5422 : begin out <= 64'b1010100011111110001001111110011100101001001010000010101100100001; end
            14'd5423 : begin out <= 64'b0010100000000100001010011100011110100101011101010010100100001101; end
            14'd5424 : begin out <= 64'b0010101110010110000101000010001010100100101100001010110000010010; end
            14'd5425 : begin out <= 64'b1010100101100100001000001010000110011010101100010010100000001111; end
            14'd5426 : begin out <= 64'b1010101001110001101000111101000100100100100110010010101010001001; end
            14'd5427 : begin out <= 64'b0010011000010010001010000001110100101000000111110010100000101000; end
            14'd5428 : begin out <= 64'b1010010010111010100110001110100000011001001000101010010011101101; end
            14'd5429 : begin out <= 64'b0010100001000010101010101000010000100001111101001010100000101011; end
            14'd5430 : begin out <= 64'b1010101110011011101011000000010010100000010101011010100101110101; end
            14'd5431 : begin out <= 64'b0010100001001010001001101100011100101001100100110010001011011011; end
            14'd5432 : begin out <= 64'b0010011011110010101010100000100000101001001111110010011010001110; end
            14'd5433 : begin out <= 64'b0010101011011000100110101000100110101011000110011010101000000111; end
            14'd5434 : begin out <= 64'b0010101111011001001001001101011000100111110111000010011101101011; end
            14'd5435 : begin out <= 64'b0010100000000000101001001110011110101010100000011010101111011000; end
            14'd5436 : begin out <= 64'b0010011011011111001010101011000010101000111111001010100101001100; end
            14'd5437 : begin out <= 64'b0010010000100100101010001111010010010100111000010010100100001111; end
            14'd5438 : begin out <= 64'b1010100110100000000111000011010010101001010101010010000110110110; end
            14'd5439 : begin out <= 64'b1010010110001001101000010100111110100100101111111010100101101100; end
            14'd5440 : begin out <= 64'b0010101001010100001010110110111100100001001110000010101101111111; end
            14'd5441 : begin out <= 64'b0010100111100111101001011111111010101011011010111010001101010100; end
            14'd5442 : begin out <= 64'b0010100011001000101010101110110000101011101010111010101010101001; end
            14'd5443 : begin out <= 64'b0010101101111000001010101011100010101011110011001010010001101110; end
            14'd5444 : begin out <= 64'b0010011101011111001001010001101110101010001110111010010101101100; end
            14'd5445 : begin out <= 64'b1010100000000110000111001011001000101010101010000010100000001111; end
            14'd5446 : begin out <= 64'b1010001001001101100111110000100110101010011101111010010000101111; end
            14'd5447 : begin out <= 64'b1010011100000100101010101101100000101010100010001010100100110010; end
            14'd5448 : begin out <= 64'b0010100001010100001010100010000110011111101000010010101111001111; end
            14'd5449 : begin out <= 64'b0010011110011100001001010000100000101000010111101010101101010010; end
            14'd5450 : begin out <= 64'b0010100011111001000101000000011000101000110011100010100110100010; end
            14'd5451 : begin out <= 64'b0010011100010101101001111100011110101010101011000010000111011111; end
            14'd5452 : begin out <= 64'b1010100011110000101010101100100100011101000100011010100100111000; end
            14'd5453 : begin out <= 64'b0010101110001100001001110001101000101010110111010010001101010100; end
            14'd5454 : begin out <= 64'b0010011000001001101010011100000010101001110100111010100110110001; end
            14'd5455 : begin out <= 64'b1010100100101010001001100010001110101010110001010010001111100111; end
            14'd5456 : begin out <= 64'b1010010110000010001000100010111110100010011100101010011000100100; end
            14'd5457 : begin out <= 64'b1010101000111111101010110111011100011110111100010010011000001111; end
            14'd5458 : begin out <= 64'b1001110011101000101010110011010100100111100110100010101011011001; end
            14'd5459 : begin out <= 64'b1010000001100101100111001011001100100011010100000001111100111010; end
            14'd5460 : begin out <= 64'b0010100001011001001010111110111110101000100000011010101010000001; end
            14'd5461 : begin out <= 64'b1010101000100000001001010001101000100011110001011010101001101011; end
            14'd5462 : begin out <= 64'b0010001100110111001000110111100110101000110001010010011100111000; end
            14'd5463 : begin out <= 64'b0010101110011111101000101000001000100011100010001010000101011000; end
            14'd5464 : begin out <= 64'b1010100010001101001000001110001010100110100000000010101101001011; end
            14'd5465 : begin out <= 64'b1010001110010100001010011110100000011010100101001010101001110011; end
            14'd5466 : begin out <= 64'b1010001010000001100111110111111100101000001000110010101010011010; end
            14'd5467 : begin out <= 64'b1001100001101100101010001111101000011100111001001010100110011100; end
            14'd5468 : begin out <= 64'b0010100100111000000111011010001110100101111111111010101110111000; end
            14'd5469 : begin out <= 64'b0010000000101001001010110001110000101011111011110010000000000011; end
            14'd5470 : begin out <= 64'b0010101000010001001001110000011110100111010011001010100101101101; end
            14'd5471 : begin out <= 64'b1010101011111000101001011101010110101010010001110010101001010110; end
            14'd5472 : begin out <= 64'b0010001011111001101001111011010000101001110101111001111000110111; end
            14'd5473 : begin out <= 64'b0010100000100101101010100101001010101001101001111010101000101011; end
            14'd5474 : begin out <= 64'b0010000011000111001001100011011000101001110100101010001010111101; end
            14'd5475 : begin out <= 64'b1010101111101101101010010010101100011101110000001010010001000101; end
            14'd5476 : begin out <= 64'b1010100000110110101001011111001000100111010001101010100110001101; end
            14'd5477 : begin out <= 64'b0010100001111100001001001110001010101011110111010001111011110111; end
            14'd5478 : begin out <= 64'b1010100001100000101010001101101110100110001010110010100000011111; end
            14'd5479 : begin out <= 64'b0010101011100001101001011001010110101010110100011010011011110110; end
            14'd5480 : begin out <= 64'b0010101100010111001010101110100000100111111010111010100011101011; end
            14'd5481 : begin out <= 64'b1010011101011100101010001001011010100000100001111010001000001101; end
            14'd5482 : begin out <= 64'b1010101011010000101001101101110000100000100011110010100101010101; end
            14'd5483 : begin out <= 64'b1010101001001001000111100101010010101011011110101010010001111010; end
            14'd5484 : begin out <= 64'b0010101001101001101010011110000100100001111100100010000101100011; end
            14'd5485 : begin out <= 64'b1010010101000011101001000001110110101000100100001001101010011111; end
            14'd5486 : begin out <= 64'b1010011111110010001001110111101110101000101100000001110101001101; end
            14'd5487 : begin out <= 64'b1010100101100001101010010110010000101000111000100001100000011001; end
            14'd5488 : begin out <= 64'b1010101000101100101010000101110010011110011101010001101011011001; end
            14'd5489 : begin out <= 64'b1010101011111101101001000000110000101011100110011010100011111111; end
            14'd5490 : begin out <= 64'b1010100101111100101001110100101010100001111000111001111000001111; end
            14'd5491 : begin out <= 64'b1010011110110110001001000001110000100011000001101010000100110101; end
            14'd5492 : begin out <= 64'b0010101110100011001010100110010010101000101010001010000110100000; end
            14'd5493 : begin out <= 64'b1010100101001001001001110101000100101000001101111010011010110011; end
            14'd5494 : begin out <= 64'b1010101000100010101001010111101000100101110100010010011011011110; end
            14'd5495 : begin out <= 64'b0010100011101011001001011001111100100000100001100010011110001110; end
            14'd5496 : begin out <= 64'b1010100000110101101000000111010100101010011111011010101011001110; end
            14'd5497 : begin out <= 64'b0010011110100110101010010110001110101011111110111010000101010110; end
            14'd5498 : begin out <= 64'b1010100100110000101001100001101000100110011001101001000110101000; end
            14'd5499 : begin out <= 64'b1010100010001010101010011000011100101001111000101010100010000010; end
            14'd5500 : begin out <= 64'b1010001100100111101001011011110100011101010000110010101111011110; end
            14'd5501 : begin out <= 64'b1001101000101111001001000000011110101011001111110010100011000010; end
            14'd5502 : begin out <= 64'b1010100111000000101000111100110000100101001000010010010101001101; end
            14'd5503 : begin out <= 64'b0010010000011110001010101100010000100110110001101010100111101000; end
            14'd5504 : begin out <= 64'b1010010010010100001010100011000000011011001001000010101110110000; end
            14'd5505 : begin out <= 64'b0010101100011011001001011110010000100101001110101010101101110001; end
            14'd5506 : begin out <= 64'b0010101010111011001010101111100000100111001111001010011110001110; end
            14'd5507 : begin out <= 64'b1001001001101010001011000111000000101011000011111010100010010101; end
            14'd5508 : begin out <= 64'b1010101111000110001001011111001100100011101000100010101100111101; end
            14'd5509 : begin out <= 64'b1010011110010010101010101000111110101001000110110010100110110000; end
            14'd5510 : begin out <= 64'b1010101010100111001010111110010000101011110001011010100010101011; end
            14'd5511 : begin out <= 64'b0010101100000111001001111000010010011101010110010010011110010111; end
            14'd5512 : begin out <= 64'b1010100100010111001010001110000100011011111011101010010011010011; end
            14'd5513 : begin out <= 64'b0001011000000101001010100101001010101001010000010010101010101111; end
            14'd5514 : begin out <= 64'b0010010001011000101000010000101100100101000001111010101010011000; end
            14'd5515 : begin out <= 64'b1010001000001001101010111101001010100001010110001010101100110011; end
            14'd5516 : begin out <= 64'b0010101001101110101010111101010100100011001011110001011001011010; end
            14'd5517 : begin out <= 64'b1010100101000110101010110101001110100011001110001010011101101100; end
            14'd5518 : begin out <= 64'b1000110100100011101010111011100110011001001100110010100011011011; end
            14'd5519 : begin out <= 64'b1000111000011100101010001010100000100111110011001001101101101001; end
            14'd5520 : begin out <= 64'b0010011101110001001010101111100000100010000101111010001000110010; end
            14'd5521 : begin out <= 64'b0010010111100100001001010011010110101011011101101010101001001001; end
            14'd5522 : begin out <= 64'b0010101010111010101001100011111000100100000001101001010010110011; end
            14'd5523 : begin out <= 64'b1010101111001110001001101000100000100110101111111010100010100111; end
            14'd5524 : begin out <= 64'b0001110111111011001000010001011010100110000101101010010011110110; end
            14'd5525 : begin out <= 64'b0010011011011011100111011000000110100001100110111001111110000101; end
            14'd5526 : begin out <= 64'b1001111001000101001010111010111010101100000010101010101001100110; end
            14'd5527 : begin out <= 64'b0010010100010101101010010101010100011101110011010010100111011011; end
            14'd5528 : begin out <= 64'b0010101000100001001000011100111100100011111100111010010111011001; end
            14'd5529 : begin out <= 64'b1010000110101110100111001000111000101010111010111010010100000101; end
            14'd5530 : begin out <= 64'b1010010010110111001010101101100100100111010001010010101011110011; end
            14'd5531 : begin out <= 64'b0010011000001100001010110000110110101000100001010010100101010101; end
            14'd5532 : begin out <= 64'b1010011101111111101000011011110110100110100110010010100111010111; end
            14'd5533 : begin out <= 64'b0010101111100001000100111110010110100101100100101010100011001010; end
            14'd5534 : begin out <= 64'b1010110000001001001010001000110110011100011001010010001000100011; end
            14'd5535 : begin out <= 64'b1010101101111000001001011000101010101011100010010010100000101111; end
            14'd5536 : begin out <= 64'b1010101000101010001010001101010100011110111110010010010101100011; end
            14'd5537 : begin out <= 64'b0010010011011011101010011101010100100110000101101010100011000101; end
            14'd5538 : begin out <= 64'b0010011110111011001000110110011000100100001100011010010000010010; end
            14'd5539 : begin out <= 64'b1010101100101000000110011001011110100101011000101010101001111110; end
            14'd5540 : begin out <= 64'b1010011100000110100111110001000010011111010110001010100000101001; end
            14'd5541 : begin out <= 64'b1010011010001000100110011111100000011110101010000010100100101000; end
            14'd5542 : begin out <= 64'b0010100111101110101010010011111100100010111100001010100101011101; end
            14'd5543 : begin out <= 64'b1010100101100111001001010001000010100001000000100010001100000010; end
            14'd5544 : begin out <= 64'b0010100101001001001001110011011010100111100100111010100010110111; end
            14'd5545 : begin out <= 64'b1010101000100010101010000010010010100100000001111010011010011100; end
            14'd5546 : begin out <= 64'b1010101111101001101001101011110010100110001101011010001101010011; end
            14'd5547 : begin out <= 64'b0010101011000000001001100101111100100001101011000010010100110110; end
            14'd5548 : begin out <= 64'b1010011110100110101010110110111000101011100110100010100100111110; end
            14'd5549 : begin out <= 64'b1010101110010000101010011010111010100101011001100010000110110010; end
            14'd5550 : begin out <= 64'b0010101101001000001010000001011100101001000100110010011100001000; end
            14'd5551 : begin out <= 64'b1010010101000111101001011100101100101001111111110010001000101101; end
            14'd5552 : begin out <= 64'b1010100101010011101010001110101010100110111110000001110100010011; end
            14'd5553 : begin out <= 64'b1010010000110111001010110001100010101001101111100010101000110011; end
            14'd5554 : begin out <= 64'b0010010010011100001010001001101000101000011110010010010101001001; end
            14'd5555 : begin out <= 64'b1010100011111111001010101100110100101010011111101010101101101111; end
            14'd5556 : begin out <= 64'b1010100000011011001010001000011110100100011000000010100111101001; end
            14'd5557 : begin out <= 64'b0010101000100111000111000101110000100000001001000010100010011100; end
            14'd5558 : begin out <= 64'b0010011000111100101010010110011010100111110110110010011111001110; end
            14'd5559 : begin out <= 64'b0010001100001100001000011101100110101010100010111010110000000001; end
            14'd5560 : begin out <= 64'b0010101111011110101010101010101010101010011001000001110111101101; end
            14'd5561 : begin out <= 64'b1001110100011010101001101110000010101011110001010010100101101101; end
            14'd5562 : begin out <= 64'b1001110100011010001001101001101100101001100000100010101000110101; end
            14'd5563 : begin out <= 64'b1001011001000111001010111001011010101011101110110010100011110101; end
            14'd5564 : begin out <= 64'b1010001001001101101010100000001010101000101001110010101001001001; end
            14'd5565 : begin out <= 64'b1010101100110101001010011101111000101001010111101010100101101000; end
            14'd5566 : begin out <= 64'b1010011011011111001010001100101110011101010111100010011110000011; end
            14'd5567 : begin out <= 64'b0010101011000100001010000101111100101010100001101010101100101101; end
            14'd5568 : begin out <= 64'b0010100110110111001001001011101000101011000111011010000010001110; end
            14'd5569 : begin out <= 64'b0010101111000001001010010100011100101001111011000010010001100110; end
            14'd5570 : begin out <= 64'b1010011001101010101000111111011100011011000101001010000011010110; end
            14'd5571 : begin out <= 64'b1010001111101001101001001110000100100101001001011010011111010011; end
            14'd5572 : begin out <= 64'b1001010010110000001010000101000100101001000011011010101101110111; end
            14'd5573 : begin out <= 64'b1010011100111000101001111010100110101100000001110010001111001011; end
            14'd5574 : begin out <= 64'b0010100010100110001010010010110000011101100000111010101011001101; end
            14'd5575 : begin out <= 64'b1010010110101100101010110010000110101011110001011010100111001000; end
            14'd5576 : begin out <= 64'b1010101100101110101010101110100110101011101001010010011110110000; end
            14'd5577 : begin out <= 64'b0001100101010110001001101010000100101000100101110010011101001111; end
            14'd5578 : begin out <= 64'b1001110100000111001010100001110000101010101001001010100100001010; end
            14'd5579 : begin out <= 64'b0010100110110101101010100111101110100111100011000010010100011110; end
            14'd5580 : begin out <= 64'b0010101110110100101010101100001000100101011111101010011000001001; end
            14'd5581 : begin out <= 64'b1010011100000101101001010001100100011110001111110001111101111001; end
            14'd5582 : begin out <= 64'b1010101000000100101010111101010000101000001000110010101000011101; end
            14'd5583 : begin out <= 64'b0010010110010110101001100010000110101010000110110001111110011111; end
            14'd5584 : begin out <= 64'b1010101011000101101000000010110110101000111010000010100101111111; end
            14'd5585 : begin out <= 64'b0010101110001101101010000111000100100100010010101010101011001010; end
            14'd5586 : begin out <= 64'b0010011101100101000111001001001110100010000101111010001011001110; end
            14'd5587 : begin out <= 64'b0010010010110101101000010100010110100100000100110010100010111111; end
            14'd5588 : begin out <= 64'b1010000111110100101001000001010110100101100111011001101111001010; end
            14'd5589 : begin out <= 64'b0010011000001101101010100000000000101011111110100010101110001100; end
            14'd5590 : begin out <= 64'b0010101100010101101001111011000000101010001010110010100010011110; end
            14'd5591 : begin out <= 64'b0010100101000101001000111011000110101001000010001010100001101000; end
            14'd5592 : begin out <= 64'b0010101101001100001010000001000000100001011100011010101110011000; end
            14'd5593 : begin out <= 64'b1010100110010010101010001100010100101000011010100010101000100011; end
            14'd5594 : begin out <= 64'b1010101011011100101010011011101100101000100111000010010010101011; end
            14'd5595 : begin out <= 64'b0001011010001110101001101000010100100100111000010010101010011010; end
            14'd5596 : begin out <= 64'b1010000100010101101010010100111000101001011101110001001001110001; end
            14'd5597 : begin out <= 64'b1010000000110101001001000100100110101000001010101010100011111011; end
            14'd5598 : begin out <= 64'b0010101101100111001010001111100100100110110010011010001100101100; end
            14'd5599 : begin out <= 64'b1010010010011100001010001111100000101011000010010010001100100001; end
            14'd5600 : begin out <= 64'b0010101010111100001010000110110100101010000100101010100000001110; end
            14'd5601 : begin out <= 64'b0001110010110010101001001011101000100111010000001010100110111010; end
            14'd5602 : begin out <= 64'b1010010010101100000111100011000110100100000001001010100000100000; end
            14'd5603 : begin out <= 64'b0010100011110010101010011110011110101000100111001010100011111100; end
            14'd5604 : begin out <= 64'b0010000011011011001010100010001100101011110101000010001011101011; end
            14'd5605 : begin out <= 64'b0010101110111010001001000001011100010110011100100010010110111001; end
            14'd5606 : begin out <= 64'b1010101000110001101010101100101000100101010110100010101011001001; end
            14'd5607 : begin out <= 64'b0010100101101110001010101000000100100001100011010010100011111001; end
            14'd5608 : begin out <= 64'b1010100001100011001001011000101110100111000100111010010001111000; end
            14'd5609 : begin out <= 64'b0010011010100101101000001110101000100101101101010010011011001000; end
            14'd5610 : begin out <= 64'b0010100110010011001010101100001100101000000001010010100010101000; end
            14'd5611 : begin out <= 64'b1010011111111001001001000000011000101000010011010010011011001110; end
            14'd5612 : begin out <= 64'b0001110111011110001010000111000110101000001110101010001111001100; end
            14'd5613 : begin out <= 64'b1010101010110001101010100000011000100110111001101010100100011100; end
            14'd5614 : begin out <= 64'b1010101011001010101010101101100110100101111010110010100101110110; end
            14'd5615 : begin out <= 64'b0010101100111010101001110001001010100110100110101010011110001000; end
            14'd5616 : begin out <= 64'b0010101010110011101001011001001110010010000001110010101100111001; end
            14'd5617 : begin out <= 64'b1010101110110110001001001011100110101011111011011001111001010100; end
            14'd5618 : begin out <= 64'b0001110010001011101010000001001000100000001010100010010010110101; end
            14'd5619 : begin out <= 64'b1010100101110001001000101001010110100110011000001010101100101111; end
            14'd5620 : begin out <= 64'b0010100101111000001010101111101110100100111100001010011011111110; end
            14'd5621 : begin out <= 64'b0010101010110110101000010011011100100000000001010010100001101000; end
            14'd5622 : begin out <= 64'b0010010000001110001001010100001010100000101110010010101011110101; end
            14'd5623 : begin out <= 64'b0010101101100111001010110010011100101010101010000010101000001010; end
            14'd5624 : begin out <= 64'b1000110001111110101010000000111000100100100111110010100001000010; end
            14'd5625 : begin out <= 64'b1010101110101100001010110110001110100000101111000010011001101010; end
            14'd5626 : begin out <= 64'b1010011011110110001010101100001000101001101010101010010001100010; end
            14'd5627 : begin out <= 64'b0010011000111011001011000000000100101010011011110010011111111100; end
            14'd5628 : begin out <= 64'b1010101001011011101010010011101100101010110111001010100101000000; end
            14'd5629 : begin out <= 64'b1010101100010010001000001010010110100111110110010010010001100000; end
            14'd5630 : begin out <= 64'b1010101111001110001010011100100100011101111101011010100100100001; end
            14'd5631 : begin out <= 64'b1010010111000110001011000000001010100111111001111001110011001011; end
            14'd5632 : begin out <= 64'b1010011110100010101010011000001110101010110111110010010010110101; end
            14'd5633 : begin out <= 64'b0010101011100001001010110000100010100000011100001010100111100011; end
            14'd5634 : begin out <= 64'b0001101001111000101010110010101100101001101011111010000000000110; end
            14'd5635 : begin out <= 64'b1010011110100000001010100010101100100111111000101010100011000001; end
            14'd5636 : begin out <= 64'b0010011111000100100110001011011100100111000101110010100101010101; end
            14'd5637 : begin out <= 64'b0010000000010010000110011101001010100001111101101010010000001001; end
            14'd5638 : begin out <= 64'b0010101010101110101001111011010110101000011111100010000100110110; end
            14'd5639 : begin out <= 64'b0010100000110111001010100101000100101010100111011010101010110100; end
            14'd5640 : begin out <= 64'b0010100111000110100110010110000000101011011110000001100110100001; end
            14'd5641 : begin out <= 64'b1010100000000001000101111110110110100101111001100010100011110110; end
            14'd5642 : begin out <= 64'b1010001111011001001010100111101000101001111000001010100101001011; end
            14'd5643 : begin out <= 64'b0010101110000001100110010010000010011110001000100000100100001101; end
            14'd5644 : begin out <= 64'b1010100101001100000111011111010110101000101011000001011100011100; end
            14'd5645 : begin out <= 64'b1010010111001010001001001011010010101001010100111010010010010110; end
            14'd5646 : begin out <= 64'b0010000101010000001010011011011010101010101110111010100010000000; end
            14'd5647 : begin out <= 64'b1010100111111110001001100110101000101001111000100010000111010100; end
            14'd5648 : begin out <= 64'b1010001100000001001001101111100100101010101100001010101010011010; end
            14'd5649 : begin out <= 64'b0010001110010110001001111001101010101010101100100010011000111100; end
            14'd5650 : begin out <= 64'b1010100010001001101001011011110110101000011101010010010001011000; end
            14'd5651 : begin out <= 64'b1010100010001111001010010101100110100111111011110010100011100011; end
            14'd5652 : begin out <= 64'b1010100000100001100110000110111000011000110110001010100000000100; end
            14'd5653 : begin out <= 64'b0010000011001000101000000010001110100100101001110010100110010111; end
            14'd5654 : begin out <= 64'b0001101111101000101010110001101000101001111100000010010000011110; end
            14'd5655 : begin out <= 64'b0010100110001000001000010000111000101011101100111010101011010000; end
            14'd5656 : begin out <= 64'b1010101000101110001000111100100100101000011111111010101001110010; end
            14'd5657 : begin out <= 64'b0010101010101101101001011000001110101010010011001010011111111100; end
            14'd5658 : begin out <= 64'b0010011100010100001010111000101010100110010100011010100110000000; end
            14'd5659 : begin out <= 64'b0010011000110001001001001110101100100100000011011010100010001110; end
            14'd5660 : begin out <= 64'b0001111110011100101010011000101000011111100101000010100011011101; end
            14'd5661 : begin out <= 64'b1010101111100000001001010111110000101011110011010010011111010000; end
            14'd5662 : begin out <= 64'b0010100101100100101010011000011110011100110010110010101001001100; end
            14'd5663 : begin out <= 64'b1010101111111001001001111011111100100101101100101010001110001101; end
            14'd5664 : begin out <= 64'b1010101000000101101010010101010110100000010000010001100000111101; end
            14'd5665 : begin out <= 64'b1010100110111010001001110100001110101011001110110010011000001100; end
            14'd5666 : begin out <= 64'b0010101011111001100111010110111100100111110111011010000010110001; end
            14'd5667 : begin out <= 64'b0010100010101110001010010111000100100001100001000010001001001110; end
            14'd5668 : begin out <= 64'b1010101010010000100111101000011010101010001111000010101101011000; end
            14'd5669 : begin out <= 64'b1010101101001100101010111001011000100101001110111001110110100010; end
            14'd5670 : begin out <= 64'b0010101000101111101010011000011110010111000001010010100011010111; end
            14'd5671 : begin out <= 64'b0010101110010111101010000000001010101010011111001010011010011110; end
            14'd5672 : begin out <= 64'b1010101110001000001010110010100110100111010000111010000011100000; end
            14'd5673 : begin out <= 64'b1010000011001010101010000011000100100111010001111010101011001100; end
            14'd5674 : begin out <= 64'b1010100000101101001010101011001110101000101110000010100011011000; end
            14'd5675 : begin out <= 64'b0010100011110101101001001000010100101000011111111010010100110000; end
            14'd5676 : begin out <= 64'b1010100110111110001001111010010110101010101101110010010011001111; end
            14'd5677 : begin out <= 64'b1010000111011100101000010010010100101011111001011010100100010101; end
            14'd5678 : begin out <= 64'b1010101000001000001010100010111110101001011010111010101010000001; end
            14'd5679 : begin out <= 64'b1010010001111011001011000100010110010000110101011010101111101111; end
            14'd5680 : begin out <= 64'b0010101000010000001010101001000100101011000011110010100100010000; end
            14'd5681 : begin out <= 64'b1010100100000001001010110011100110101011101010110010001000110100; end
            14'd5682 : begin out <= 64'b0010101110110010101001101001101000101011011001101010000101110100; end
            14'd5683 : begin out <= 64'b0010000010001100101010101101011110101000011010011010001111111000; end
            14'd5684 : begin out <= 64'b1010000011001010101010000111100000101001110000011010100011010011; end
            14'd5685 : begin out <= 64'b0010010010111000101010110101100010011111001101100001110101100110; end
            14'd5686 : begin out <= 64'b0010010001111110101010011011101100101011011111101010101011010001; end
            14'd5687 : begin out <= 64'b0010011000101000001010101111011010101011011000100010010110010010; end
            14'd5688 : begin out <= 64'b0010100010111001100111011100111110101001001100100010100101010110; end
            14'd5689 : begin out <= 64'b0010010111101011101001000110111010001010000001011010010000000000; end
            14'd5690 : begin out <= 64'b0010101011100110001001001101111110101001101111110010000011010011; end
            14'd5691 : begin out <= 64'b0010001101100001100101111110111010100100010110011010101111010111; end
            14'd5692 : begin out <= 64'b1010000010101110001010101010101010101000010101100010010011011010; end
            14'd5693 : begin out <= 64'b0010010010101111101010111101000010100101011110010001110110101101; end
            14'd5694 : begin out <= 64'b1010101010000110101010111101000000011011011110011010101110010110; end
            14'd5695 : begin out <= 64'b0010100111100000101000010110001100011010000110001001101001100010; end
            14'd5696 : begin out <= 64'b1010100000011110101001001011100100100001001011101001100000001000; end
            14'd5697 : begin out <= 64'b0010101101000110101001101110010010101011110001000010010110110101; end
            14'd5698 : begin out <= 64'b0010100001011111001010001100101110101100000000001010001101011110; end
            14'd5699 : begin out <= 64'b0010010001101110101001000101100010101010100011100010010010000100; end
            14'd5700 : begin out <= 64'b1010010111000001101010000001000110011000110011100010010101110110; end
            14'd5701 : begin out <= 64'b1010100001001101000111111001111100101001011001100010010100000111; end
            14'd5702 : begin out <= 64'b0010000001101011101010111011111010100110101011001010100010001001; end
            14'd5703 : begin out <= 64'b0001101010110000101010100000010110101010011110110010101000000000; end
            14'd5704 : begin out <= 64'b1010101011001111101001111010101110100110001001010010100111110101; end
            14'd5705 : begin out <= 64'b1001100010010110101001011111101010101001011011000010011010000010; end
            14'd5706 : begin out <= 64'b1010101110001011001001101001010000100001100001100010011011010011; end
            14'd5707 : begin out <= 64'b0010100010101100001010110000111010101001010111111010001010010011; end
            14'd5708 : begin out <= 64'b1010101111010110001010000000111100101000110100100010011001110010; end
            14'd5709 : begin out <= 64'b0010100010010010001010110010101100100110000110010010100100111000; end
            14'd5710 : begin out <= 64'b1010100110000000001000110110111110011000011001111010100100011110; end
            14'd5711 : begin out <= 64'b1010000111010011101010011011011010011110001111110010100111010101; end
            14'd5712 : begin out <= 64'b1010100110000111001001100111101000011100111001000001100101001111; end
            14'd5713 : begin out <= 64'b0010100000001111001010000011001110100110100010111010100001101101; end
            14'd5714 : begin out <= 64'b0010000011001010101000100101000110101001111111001010100101011101; end
            14'd5715 : begin out <= 64'b0010101111100000000110000110110110101001110011000001110100011111; end
            14'd5716 : begin out <= 64'b0010011011001001101000011100011100101001101001010010100110100111; end
            14'd5717 : begin out <= 64'b1001101101001101101010101000000100101000100100110010101011111000; end
            14'd5718 : begin out <= 64'b1010000000100001001010101100100000100100011111001010010010101010; end
            14'd5719 : begin out <= 64'b0010001010110001101001110001100100011000011011001010100011100100; end
            14'd5720 : begin out <= 64'b0010100110010110001000001111011100101001010000010010010111101111; end
            14'd5721 : begin out <= 64'b1010011010011010001011000001111000101001011101110001110001000110; end
            14'd5722 : begin out <= 64'b1010100111101001000111010101100110100000000000101010011111101000; end
            14'd5723 : begin out <= 64'b0010101111000111101000000100100100100010000001000010000001110001; end
            14'd5724 : begin out <= 64'b1010101110111100001010110110001110100101000110101010101101000110; end
            14'd5725 : begin out <= 64'b0010101100000010100111101110110110100000111001101010100011110001; end
            14'd5726 : begin out <= 64'b0000000101111110101001011111011010100010010010101010101000011001; end
            14'd5727 : begin out <= 64'b0010100001111111001010101101000110101011110101000010010011101011; end
            14'd5728 : begin out <= 64'b1010011011110010001010001011000100101011010110100010011000000011; end
            14'd5729 : begin out <= 64'b1010011111101000001010100100000000000010000101101001111001101110; end
            14'd5730 : begin out <= 64'b1010100000101010101001001110111110101010010111111010010110010100; end
            14'd5731 : begin out <= 64'b0010100110110111000111000010110000101011100000111010100100110001; end
            14'd5732 : begin out <= 64'b1010101001110011001001110100000110100011101101010001010110001111; end
            14'd5733 : begin out <= 64'b1010101010010111001010110001011000101001011010000010010010000001; end
            14'd5734 : begin out <= 64'b0010101110001101101001101010001110101000110001100010010111001111; end
            14'd5735 : begin out <= 64'b1010101100000000101001110111001110100010010001010010100011000010; end
            14'd5736 : begin out <= 64'b1010000010011111001001111010101100101010001001011010100101001011; end
            14'd5737 : begin out <= 64'b1010010010000011101010100110001010101011011010100010101110111110; end
            14'd5738 : begin out <= 64'b1010011100010111000111010111111010010001000111010010100110110111; end
            14'd5739 : begin out <= 64'b1010011000101000101001011101110000101010000011011010001100011001; end
            14'd5740 : begin out <= 64'b0010100001001111100100011010110000100100100010101010000100110110; end
            14'd5741 : begin out <= 64'b1010101100101001001010100011111010100101101011100010010010101010; end
            14'd5742 : begin out <= 64'b0000011110011110101010100010011010100100101100001010100001101011; end
            14'd5743 : begin out <= 64'b0001101101001100001010100001001010100111010011000010100101010101; end
            14'd5744 : begin out <= 64'b1010001110111001101010100100111100101001011001100010011101101100; end
            14'd5745 : begin out <= 64'b1010100111111100001010100101000010100010101101111010101111110101; end
            14'd5746 : begin out <= 64'b0010000000011010101001101100100110101011101000101010101101001111; end
            14'd5747 : begin out <= 64'b1010001010100000101000101011101000100101110111010010001110111101; end
            14'd5748 : begin out <= 64'b0010000110100011100110100011010000101000000111111010101101001000; end
            14'd5749 : begin out <= 64'b1010101111111000001001101001011110010111011001110010100101100101; end
            14'd5750 : begin out <= 64'b0010101000111010101001010010000110101001000110101010101000110101; end
            14'd5751 : begin out <= 64'b1010100001001010100111011101011110100110001110111010101111000101; end
            14'd5752 : begin out <= 64'b1010010101110010101010100111111000101001010110101010010000000111; end
            14'd5753 : begin out <= 64'b0010100101010100001001110000110000101010100001001010101111001011; end
            14'd5754 : begin out <= 64'b0010101001101000101010110011110100101010111010010010001110100100; end
            14'd5755 : begin out <= 64'b1010011101001100001000100001101110101000111111010010100100110100; end
            14'd5756 : begin out <= 64'b0010101011010111101001101100001100101000001110001010101000010010; end
            14'd5757 : begin out <= 64'b1010100011111001101010001101010110101010110001011010000000001100; end
            14'd5758 : begin out <= 64'b0010101001110111001010101000011010100101000001101001110000011001; end
            14'd5759 : begin out <= 64'b1010000010001100101010100110011110011111011111100010000110101111; end
            14'd5760 : begin out <= 64'b0010101111111000101001010111100000010101011111001010011000111000; end
            14'd5761 : begin out <= 64'b1010100100011001001010010000101100101001101011100010100001110101; end
            14'd5762 : begin out <= 64'b0001100001101011001010101101000000001111011000001010010000010101; end
            14'd5763 : begin out <= 64'b1010100010101111001011000011001110011001000001111010101000011011; end
            14'd5764 : begin out <= 64'b0010010000100001001010101111000110101011001010100010000000011001; end
            14'd5765 : begin out <= 64'b1010101111010111101010011101111010100010011110100010101100001111; end
            14'd5766 : begin out <= 64'b1010101010100010001001100111110100101000010011100010100011110100; end
            14'd5767 : begin out <= 64'b1010100011110011001010101001001010100100110101011010011101010000; end
            14'd5768 : begin out <= 64'b1001110110001010101001101001110010100110100100000010001000001000; end
            14'd5769 : begin out <= 64'b0010100110010100001000100011000010011100110111100010101100100011; end
            14'd5770 : begin out <= 64'b1010100111110001101010001100100010101011111111111010101011001000; end
            14'd5771 : begin out <= 64'b1010011010101101001001011101000100101000001011111010101100001110; end
            14'd5772 : begin out <= 64'b0010101010110101001010100110110110101001000110110010011001101110; end
            14'd5773 : begin out <= 64'b1010011010011111100110000110111110101001011100100010011111000011; end
            14'd5774 : begin out <= 64'b1010100100010000000101111011001100100000011110001010100001110101; end
            14'd5775 : begin out <= 64'b0010011110111011101010110101111110100001001011001010010110100101; end
            14'd5776 : begin out <= 64'b1010010100100101101010101100100000100111110100001010100111110000; end
            14'd5777 : begin out <= 64'b0010010101001101001010100100011110101011110010001010100110100000; end
            14'd5778 : begin out <= 64'b1010101111111011000100110110100000101010110010010010100110010000; end
            14'd5779 : begin out <= 64'b0010101000001110101010111000101000100000101011010010010001101110; end
            14'd5780 : begin out <= 64'b0010011100110111001010011011010000100001010101011010100110000111; end
            14'd5781 : begin out <= 64'b0010101011001110101010101001101000100111111111001010010100001001; end
            14'd5782 : begin out <= 64'b0010101110100000000111100100011110100101010101010010100110001101; end
            14'd5783 : begin out <= 64'b0010101011100100001010000111000100100011001100111010011101010010; end
            14'd5784 : begin out <= 64'b0010101011001000000111101111100100101010110110101010000110001100; end
            14'd5785 : begin out <= 64'b1010010101100000001010110101100000101000001100001010010101111001; end
            14'd5786 : begin out <= 64'b1010100100010000101010101001111010100101011000111010100111110101; end
            14'd5787 : begin out <= 64'b1010100000010101001000000100000100100001100100110010100001110101; end
            14'd5788 : begin out <= 64'b0001100001110110001010000110101010101001001111111010000100000011; end
            14'd5789 : begin out <= 64'b1010101001100001101010000101111010101000001101011010001111100101; end
            14'd5790 : begin out <= 64'b1001101001100110101010001001000000101001111010110010101111011110; end
            14'd5791 : begin out <= 64'b1000100001101000001001101010110100100011111111111001110101101011; end
            14'd5792 : begin out <= 64'b1010100000011101001001010110011010101010111011101010010000100001; end
            14'd5793 : begin out <= 64'b1010100100110101001010100010101000100100100010100010100000101010; end
            14'd5794 : begin out <= 64'b1010011010100000101010110111001100100110001011000010101110101001; end
            14'd5795 : begin out <= 64'b0010100100101101001010011010001000100110100111110010100100101000; end
            14'd5796 : begin out <= 64'b0010011111011010001000001011101000100000001011010010001110000000; end
            14'd5797 : begin out <= 64'b0001111111001101101010010010010010101011111111111010101010010011; end
            14'd5798 : begin out <= 64'b0001111000010001001001111000010010101000010000011010101000011001; end
            14'd5799 : begin out <= 64'b0010100110011001101010111111110110100110000111001010101001111100; end
            14'd5800 : begin out <= 64'b1010011100100110000101000001000010101001101010100010000001010001; end
            14'd5801 : begin out <= 64'b0010100001111001001001110001101000101000011101100010101000011101; end
            14'd5802 : begin out <= 64'b1010100110001000001010111110011000101000110010010010101001100010; end
            14'd5803 : begin out <= 64'b1010101100100001101010110101100110101010000000100010101000000001; end
            14'd5804 : begin out <= 64'b1010011110011100001000111010110110101000101111010010011000010001; end
            14'd5805 : begin out <= 64'b0010100110010101000111111110000100101010000100000010011011100101; end
            14'd5806 : begin out <= 64'b0001011011000001101000101100010100101000110101100010011101110111; end
            14'd5807 : begin out <= 64'b1010011101100110001010000100110100001100010100010010000011111100; end
            14'd5808 : begin out <= 64'b0010010111100101101001111111001100100011111100001010010101111001; end
            14'd5809 : begin out <= 64'b0010001011110000001001001001101100100100001000110010101010100001; end
            14'd5810 : begin out <= 64'b1010100000100011001010010000010000101010011111010010100011110111; end
            14'd5811 : begin out <= 64'b0010011000111100000111000110011110101000001101110010011110100011; end
            14'd5812 : begin out <= 64'b0010101111000111001001011001011000100110110001001010011010101110; end
            14'd5813 : begin out <= 64'b1010010000011011100111001110110100100100001110000010000110011011; end
            14'd5814 : begin out <= 64'b1010000111101111001000001101011010101001101110011001100011010101; end
            14'd5815 : begin out <= 64'b0010101110000110101010100110100000100111010010100010100011011000; end
            14'd5816 : begin out <= 64'b1010010100010101001001110111010000101000110100000010011001111001; end
            14'd5817 : begin out <= 64'b0010010011000001101001101101110010100111001110010010101110010100; end
            14'd5818 : begin out <= 64'b0010101111011010001000101000001010101010111001111000101100001001; end
            14'd5819 : begin out <= 64'b0010101111101001001011000001100110101000111110100010010100010010; end
            14'd5820 : begin out <= 64'b1010100111100101001010111111111010101001011011101010100110001011; end
            14'd5821 : begin out <= 64'b0010010100011011101010001011000110011111111110100001100011110001; end
            14'd5822 : begin out <= 64'b1010100001111000000111111000111100010100010111111010101100100001; end
            14'd5823 : begin out <= 64'b1010010010110111001010111000101010100111111100101010001001100000; end
            14'd5824 : begin out <= 64'b1010011110100000101010100000011110100111101000101010101100111000; end
            14'd5825 : begin out <= 64'b1010100000011101101000111100000000100100000110100010010011001111; end
            14'd5826 : begin out <= 64'b0010100111101111101000101011111000101011011111101010100100101100; end
            14'd5827 : begin out <= 64'b0010101010001101000110011010001000101000011110110010100011000110; end
            14'd5828 : begin out <= 64'b0010001010111110001010101001110100101001111110001010001010100011; end
            14'd5829 : begin out <= 64'b1010011000000110000111110001000000101010101010011010011011000000; end
            14'd5830 : begin out <= 64'b1010011011101101101001010000111010100011100100000010101101111000; end
            14'd5831 : begin out <= 64'b0010010101100111001010110011111000100100010001000001100110001011; end
            14'd5832 : begin out <= 64'b1010100110110110101010101001000100101001001001000010101011110011; end
            14'd5833 : begin out <= 64'b1010101101111011001010011011100010100011101010100010101000111011; end
            14'd5834 : begin out <= 64'b0010100101000101001010010110110010101011110101010010011000110011; end
            14'd5835 : begin out <= 64'b1010101110011101001001011110110100100110101010001010101010110001; end
            14'd5836 : begin out <= 64'b1000111001100000101001000010110110100101111101100010001110101111; end
            14'd5837 : begin out <= 64'b1010001000100100001010100101100100101010100001011010101010110011; end
            14'd5838 : begin out <= 64'b0010101111110000101001011100110100100110100000101010101111111010; end
            14'd5839 : begin out <= 64'b0010100100011100001001001011101100101010011101000010100110000101; end
            14'd5840 : begin out <= 64'b0010010110100011001010111111101110101010001100000010011010111110; end
            14'd5841 : begin out <= 64'b1010011110011000101010110001110110101001000110101010001000100010; end
            14'd5842 : begin out <= 64'b0010011011010100101001101101010100100011110101011010101111011100; end
            14'd5843 : begin out <= 64'b1010010101100000101010000101100000101000110011110010101100100110; end
            14'd5844 : begin out <= 64'b0010101010100101101010000101001000011111001101111010101111010101; end
            14'd5845 : begin out <= 64'b1010100010101111100011110111010010100101111111000010011011000100; end
            14'd5846 : begin out <= 64'b1010101100001011001010001011011000100001100110111010101010110100; end
            14'd5847 : begin out <= 64'b0010100101110001101000101111101000100011111011000010010001110011; end
            14'd5848 : begin out <= 64'b1010100011101101001010001101111110011010011110100001111111011010; end
            14'd5849 : begin out <= 64'b1010101011010010001011000001100100101011111000100001111111001111; end
            14'd5850 : begin out <= 64'b1010101001001011001000100100010000011000011100111010100101000000; end
            14'd5851 : begin out <= 64'b0010010000010110101010100000101000101011111111110010001011010101; end
            14'd5852 : begin out <= 64'b0001010100011010001010101001111110100110100010010010010000100101; end
            14'd5853 : begin out <= 64'b1010101000110101001010110001101000100111110010011010101110110100; end
            14'd5854 : begin out <= 64'b0010101110101110001001000010011100100100111100111010011010111011; end
            14'd5855 : begin out <= 64'b0010101010110011001001100111011000100110001001001010101010001001; end
            14'd5856 : begin out <= 64'b0010010101100010101010110110000000100110100111110010100011101101; end
            14'd5857 : begin out <= 64'b1010100011111111101001110001001010101010001100011001110011000011; end
            14'd5858 : begin out <= 64'b1001100010000001001001110100000010101010111100011010100011110010; end
            14'd5859 : begin out <= 64'b0010010111110000101010111010101100011101111001011010000001110011; end
            14'd5860 : begin out <= 64'b1010101000110101101010001010011010101010110111010010101010101011; end
            14'd5861 : begin out <= 64'b0010001000111100101010001010001000101001110000100010101101011110; end
            14'd5862 : begin out <= 64'b1010101100000111000100011011101010101000111101100010100010011000; end
            14'd5863 : begin out <= 64'b1001111010111110001011000000111000100111101011010010000111111111; end
            14'd5864 : begin out <= 64'b0010100010001101101010000001010000101011000110001010100111011011; end
            14'd5865 : begin out <= 64'b1010101010110111001001110011110000100011011111000010011000001110; end
            14'd5866 : begin out <= 64'b0010100010101010101010101000101010100010101100001010101100000011; end
            14'd5867 : begin out <= 64'b1010010010110011001010100011001010100110111111011010011101010001; end
            14'd5868 : begin out <= 64'b1010101000111010000111001101101110101001000111011001100110000110; end
            14'd5869 : begin out <= 64'b0001110001000010001000100010101110100000001111000010001011101100; end
            14'd5870 : begin out <= 64'b0001110110110110101010100011110110101010000011010010100111100100; end
            14'd5871 : begin out <= 64'b1010000001000101001010100010010110101011110100000010101101101110; end
            14'd5872 : begin out <= 64'b0010011011010000000011100010100110100111111011010010101101010001; end
            14'd5873 : begin out <= 64'b0001101001011010101001100011111100100111000000001001101110111101; end
            14'd5874 : begin out <= 64'b1010101100110001001000010100001100101010110000000010101111110111; end
            14'd5875 : begin out <= 64'b1010101110110011101000101011010110100101101011011010011011000110; end
            14'd5876 : begin out <= 64'b1010101111110110101001001100011110100001100110100010010001011001; end
            14'd5877 : begin out <= 64'b0010101010100100001010011001111010101010100011101010101001010110; end
            14'd5878 : begin out <= 64'b0010011100000001001010010100101000101011001010011010011001100101; end
            14'd5879 : begin out <= 64'b0010100000111111001001000011111010100111011010001010101000101110; end
            14'd5880 : begin out <= 64'b1010010001010010101010010010110000011110000010100001010011010000; end
            14'd5881 : begin out <= 64'b0010101110111110100101101010111010101000001111010010101000101001; end
            14'd5882 : begin out <= 64'b0010011011000111101001011111101000101001011100110010101111001001; end
            14'd5883 : begin out <= 64'b1010101011100111001000000000011010100100100111100010101101011011; end
            14'd5884 : begin out <= 64'b1001110111011001101001110100010000101001101111100010101111010100; end
            14'd5885 : begin out <= 64'b0010101111111111100110001011100110011100001011000010001011100100; end
            14'd5886 : begin out <= 64'b1010010010010001001001101110010010100010111010100010100110010100; end
            14'd5887 : begin out <= 64'b1010101010001011100111000000011010100111001100000010010100011111; end
            14'd5888 : begin out <= 64'b1010100011100110101000000111000010101011101011011001101010110101; end
            14'd5889 : begin out <= 64'b0000001110101011001010010100100010101010110001111010100011010101; end
            14'd5890 : begin out <= 64'b1010100011010111001000110000100000100110100000001010000000101100; end
            14'd5891 : begin out <= 64'b0010010001111101001010101110011110100000101000101010101010010010; end
            14'd5892 : begin out <= 64'b1010101001101100001010110010001110101000000111010001110001101100; end
            14'd5893 : begin out <= 64'b0010011101101101101010000111110000101010000001101010001001101101; end
            14'd5894 : begin out <= 64'b0010010101110100001001100111001000101000010011110010011111111011; end
            14'd5895 : begin out <= 64'b1010010100101000101010011011100100010111110100010010010110001110; end
            14'd5896 : begin out <= 64'b1010101100110110101001000100000000101001111000010000000010001000; end
            14'd5897 : begin out <= 64'b0010010011101010101001100011111100100001111001011010010110001001; end
            14'd5898 : begin out <= 64'b0010101011001011001010101010010110100000100100010010100011001101; end
            14'd5899 : begin out <= 64'b1010000000110101001010010110000000010111101101000010001101000001; end
            14'd5900 : begin out <= 64'b1010000101111011101010000000001010100111100110111010100010110001; end
            14'd5901 : begin out <= 64'b0001101101001100101001010011010010101001110000000010010001101010; end
            14'd5902 : begin out <= 64'b1010100000011010101010100001101100100100100010000001101010011011; end
            14'd5903 : begin out <= 64'b0010101100111101001001111110100100100100100100001010011101010101; end
            14'd5904 : begin out <= 64'b0010101101110100101010101001110000101000000010101010101100001000; end
            14'd5905 : begin out <= 64'b1010101001010110101010011011111000100000000001000010101010000101; end
            14'd5906 : begin out <= 64'b0010100110110100001001110101110100100110010101110010100111101010; end
            14'd5907 : begin out <= 64'b1010000001110101001000100101111110101011111001100010010111101101; end
            14'd5908 : begin out <= 64'b0010101000111000001010000001000010100101101110101010001101010001; end
            14'd5909 : begin out <= 64'b0010100001111010101000101000111100101011100111100010101101000110; end
            14'd5910 : begin out <= 64'b1010100101010110001010001101110100100100110000001010010111110000; end
            14'd5911 : begin out <= 64'b1010011000001011100111011011111000101001101010111010100100100010; end
            14'd5912 : begin out <= 64'b1010101110110111101001011100101100100111001101101010011011000100; end
            14'd5913 : begin out <= 64'b0010101001111011101000001010100100101001011111110010011100110010; end
            14'd5914 : begin out <= 64'b0010001110101001100111001010010100101000001111011010010011111100; end
            14'd5915 : begin out <= 64'b0010011111010011101010010011001000101010110010100010011111000100; end
            14'd5916 : begin out <= 64'b0001110100001001001001111110010110101001100000011010001100011010; end
            14'd5917 : begin out <= 64'b1010100010100100101010100110000100101100000010010010101001000010; end
            14'd5918 : begin out <= 64'b1010101110011001101010010100111010101001110111101010101010111010; end
            14'd5919 : begin out <= 64'b0010101100001110000111001001101010011111110101010010101111001110; end
            14'd5920 : begin out <= 64'b0010010011101100101010101111100100101000110110010010101010001110; end
            14'd5921 : begin out <= 64'b0001111010010010001010000100111010100100000000001010010100101011; end
            14'd5922 : begin out <= 64'b1010100000001110101010111000011000100101111111111010010001001010; end
            14'd5923 : begin out <= 64'b0010011101111010101010110100110010011100001000001001111101110110; end
            14'd5924 : begin out <= 64'b1010010000010011000101000010001100101011001001100001111110101001; end
            14'd5925 : begin out <= 64'b1010001111010000101011000001000000101001100110000001101111001001; end
            14'd5926 : begin out <= 64'b1010101000100111101010110100101110011111010000000010001001110110; end
            14'd5927 : begin out <= 64'b0010101011011001001010101101100000101010000110101010010000100101; end
            14'd5928 : begin out <= 64'b1010101000011111101000110111100110101001101111011010101100100100; end
            14'd5929 : begin out <= 64'b0010100010101101001000101101110000101010010011011010001001001100; end
            14'd5930 : begin out <= 64'b0010010100000111100111010101110000100111000101010010101111001001; end
            14'd5931 : begin out <= 64'b1010001000001011001011000000001110100101001110101001111011101110; end
            14'd5932 : begin out <= 64'b0010101111100001001010001111101100011101000011011010100111110100; end
            14'd5933 : begin out <= 64'b0010001110111110001010100111001110011001001111001010100111010110; end
            14'd5934 : begin out <= 64'b1010010000110010100111101011000100101001110001000010010111111111; end
            14'd5935 : begin out <= 64'b1010011011100110101001101010101100101000110000011010101010100101; end
            14'd5936 : begin out <= 64'b1000100111010111001010100010001100101011100110010010011010011110; end
            14'd5937 : begin out <= 64'b0010101101101001101010001100000010101011011000111010101010111101; end
            14'd5938 : begin out <= 64'b0010100011011111101001010100100100101000010001110010011110010111; end
            14'd5939 : begin out <= 64'b1010100011010010101010010100110000101000110111001010100000110101; end
            14'd5940 : begin out <= 64'b1010100010101001101000110101001110011001001101001010101101111100; end
            14'd5941 : begin out <= 64'b0001011101000011101001000111010110101100000010101010000000110100; end
            14'd5942 : begin out <= 64'b1010000100111111101001010001101100101000001100001010010100000000; end
            14'd5943 : begin out <= 64'b0010101100010111101010101110010010101000111110110010000110101111; end
            14'd5944 : begin out <= 64'b1001110101011101001010000000111110100011101110000001100000011001; end
            14'd5945 : begin out <= 64'b1010101010111100101000111001001010100110110100110010101011011110; end
            14'd5946 : begin out <= 64'b1010011100100011001000110101000000101010010111011010001010110010; end
            14'd5947 : begin out <= 64'b0001110000101000001010010010100010100001100110001010011011100100; end
            14'd5948 : begin out <= 64'b1010101111011000001001111011101010100000100000011010011101101011; end
            14'd5949 : begin out <= 64'b1010100001001110101010001110100100101010110101101010011010111101; end
            14'd5950 : begin out <= 64'b1010011100110001001001000100011110101001011001111010010010011110; end
            14'd5951 : begin out <= 64'b1010001010101111001000111100010010101010101111000010011100010000; end
            14'd5952 : begin out <= 64'b0010100010111110001000011000001100101010001101111010100101010111; end
            14'd5953 : begin out <= 64'b1010000001001100001010101111000100101010101100110010010111111010; end
            14'd5954 : begin out <= 64'b0010100011101001001010111001101000101001010001110010100011010100; end
            14'd5955 : begin out <= 64'b1010001011001110001010100011110000101000001000100010000001001101; end
            14'd5956 : begin out <= 64'b1010100011011010101001000001010110100011101111001010011010011111; end
            14'd5957 : begin out <= 64'b1010100110111101001001001010110100100011110000111010001001101111; end
            14'd5958 : begin out <= 64'b0010101100110101100011100000100000101010011101011001010100111111; end
            14'd5959 : begin out <= 64'b1010101011001101001001001011111110100111001101010001110111101100; end
            14'd5960 : begin out <= 64'b0010100010100011001010011000011100101001100000110010101011001001; end
            14'd5961 : begin out <= 64'b1010100110111000101010100101011000101001101010111010001100001100; end
            14'd5962 : begin out <= 64'b1001010011101110001010000010111010101011010111000010100100000001; end
            14'd5963 : begin out <= 64'b0010010110111111000101000001000010101001110101001010100000000111; end
            14'd5964 : begin out <= 64'b1010011101001111001010110110100100101011111010110010010101100101; end
            14'd5965 : begin out <= 64'b1001111010100001001000101111110000011001111000111010100001100100; end
            14'd5966 : begin out <= 64'b0010101100111101001010101110110100101010110010010010101010110000; end
            14'd5967 : begin out <= 64'b0010011110110111101001111010110100101011101011110010101001011011; end
            14'd5968 : begin out <= 64'b1010101001001111101010011100000010100101101000110010101100000100; end
            14'd5969 : begin out <= 64'b1010011010010011001010010000011010101010001000000010010100001010; end
            14'd5970 : begin out <= 64'b1010100011111001101010010111111010101011110110000010101101000100; end
            14'd5971 : begin out <= 64'b1010010011111110101010001110100100011100001111011001111100101010; end
            14'd5972 : begin out <= 64'b1010101000011111001000001010101100100100110000101010100011001011; end
            14'd5973 : begin out <= 64'b1010100001100100001010001111110100100110010001111010010000000110; end
            14'd5974 : begin out <= 64'b1001111101011100001010110110001010101011111000011001110100111011; end
            14'd5975 : begin out <= 64'b0010000111001100001010100100111010100010100000100010011010101010; end
            14'd5976 : begin out <= 64'b0010010101000001101001100101010100101011000101100010001011100110; end
            14'd5977 : begin out <= 64'b1010101111001010101010100110011000101001111101101001101000010100; end
            14'd5978 : begin out <= 64'b1010101000010001101001001011000100101011010001111010011000100011; end
            14'd5979 : begin out <= 64'b1010010110000000101000100010110010100111101101001010011010001101; end
            14'd5980 : begin out <= 64'b0010101110000111101010110101101100100111100000010010001110011110; end
            14'd5981 : begin out <= 64'b1010100101100100001010100010110110100101000111001010100010110110; end
            14'd5982 : begin out <= 64'b0010001110011000000111100100000000101010011101101010100001010010; end
            14'd5983 : begin out <= 64'b0010101110000010101001010110110110100011010010110010110000001000; end
            14'd5984 : begin out <= 64'b0010010010000000101001100111111000100110001101010010100111011101; end
            14'd5985 : begin out <= 64'b0010010000111100101010101010110000101001100100100010101100111100; end
            14'd5986 : begin out <= 64'b1010101100110011001010101011110100011010111100011010100011010111; end
            14'd5987 : begin out <= 64'b0010101001111010101010110011111110101011000000111010000001111011; end
            14'd5988 : begin out <= 64'b0010010000011111101001000011110100010001000010110010100000101001; end
            14'd5989 : begin out <= 64'b1010100110110101001010101000000110101001101000010010011010110101; end
            14'd5990 : begin out <= 64'b0010010011010011101011000000100010011101111110001010011111001110; end
            14'd5991 : begin out <= 64'b1001111100111000101001101000010110100110000111111010001101110000; end
            14'd5992 : begin out <= 64'b1010101001010111001010100000010000101010100000001001100001001001; end
            14'd5993 : begin out <= 64'b0010011111100111001010100001100110011011100000100010011110000010; end
            14'd5994 : begin out <= 64'b0010101000100011101001000001010100101000000100110010100010110001; end
            14'd5995 : begin out <= 64'b1010100111011001001010000001001000101011001011111010100101100100; end
            14'd5996 : begin out <= 64'b0010011101001100101010110100110110101010111001101010100101011010; end
            14'd5997 : begin out <= 64'b0001101111011101100111011100101000100110110100110010100011110010; end
            14'd5998 : begin out <= 64'b1010100010001010001000010010001000100001001010100010101000010100; end
            14'd5999 : begin out <= 64'b0010011101000010101010101010110110101010000000100010100000010000; end
            14'd6000 : begin out <= 64'b0010100011000101001000011010100100100111001011101010100110100101; end
            14'd6001 : begin out <= 64'b0010101110101100001010101000101100100011001100101010100011110010; end
            14'd6002 : begin out <= 64'b0001111011001101001001111100011010100100101010101001110100101001; end
            14'd6003 : begin out <= 64'b1010011101011000101000101111010110101011101011110010101000000101; end
            14'd6004 : begin out <= 64'b0010000011111001100111100111111010100111111100011010100011101111; end
            14'd6005 : begin out <= 64'b1010101110101001001010001010110000100110000110111010100111000100; end
            14'd6006 : begin out <= 64'b1010100100110000001001000110110000100110101000001010101110010000; end
            14'd6007 : begin out <= 64'b0010100010100111101001101101110000100100111011110010100111010100; end
            14'd6008 : begin out <= 64'b0010000001010101001010110011001110100010101001110010101011110101; end
            14'd6009 : begin out <= 64'b1010100110011101101001011100010000100010010010111001110010101101; end
            14'd6010 : begin out <= 64'b0010011011101011101010000101110110010001100011110010010111000001; end
            14'd6011 : begin out <= 64'b0010100001010111101010101100111000100110100110011010100011000011; end
            14'd6012 : begin out <= 64'b1010101010001101101001011011010110101001110000110010000001101100; end
            14'd6013 : begin out <= 64'b0010011101111111000000001110011010101010111110110010100011111011; end
            14'd6014 : begin out <= 64'b1010100110000111101010110111000110011100001011011010010000011110; end
            14'd6015 : begin out <= 64'b0010011010011111001001000001011010101011110111011010101100010010; end
            14'd6016 : begin out <= 64'b0010101001001001001001001011100010100111100000111010000011011110; end
            14'd6017 : begin out <= 64'b0010100100011000001010110110001110100110010001101010010101000101; end
            14'd6018 : begin out <= 64'b1010101001111110000110110010110000101010110101010010000111001010; end
            14'd6019 : begin out <= 64'b1010101110011000000111101110001010011111111011111010010110010101; end
            14'd6020 : begin out <= 64'b0001111011001111101001000100100000100101100110010010010011000111; end
            14'd6021 : begin out <= 64'b0010110000010000101001111101001010101001100010000010010101110011; end
            14'd6022 : begin out <= 64'b1010001101000101101010100010111010101010011110101010000011001110; end
            14'd6023 : begin out <= 64'b0010100010100010101001101000001000101001101100010010011011001101; end
            14'd6024 : begin out <= 64'b0010001011010100101001001111111100101011100011000010100010000100; end
            14'd6025 : begin out <= 64'b1010100000011101100111010100100010001110101001000001101100000100; end
            14'd6026 : begin out <= 64'b1001110010001001001010000011000100100111011000011010000001001111; end
            14'd6027 : begin out <= 64'b1010011010100101101001100111001100100011010001110010010001011100; end
            14'd6028 : begin out <= 64'b0010001101110101001010100010111000100111001000101010101100011001; end
            14'd6029 : begin out <= 64'b0010101000101001101010110101100000100011101001000010100000111010; end
            14'd6030 : begin out <= 64'b1010100011100010000111110011101110101000110101011010000101110010; end
            14'd6031 : begin out <= 64'b1010011111101111101010111101110010101000000001010010101110000111; end
            14'd6032 : begin out <= 64'b1010100111100000001000101110101110101100000011110001110010101110; end
            14'd6033 : begin out <= 64'b1010101101011010100111101111100110101001000111101010101011110101; end
            14'd6034 : begin out <= 64'b0010100100010000100111110011111110101001011110111010100010101001; end
            14'd6035 : begin out <= 64'b1001111000111001001000010101110000101001010001101010011010011100; end
            14'd6036 : begin out <= 64'b0010100101110011001010111101101010101011011010001010100000101111; end
            14'd6037 : begin out <= 64'b0010101100111100101010000000111010011111010100100010011111000110; end
            14'd6038 : begin out <= 64'b0010100001110111101000100111111010101001011000011010101001000010; end
            14'd6039 : begin out <= 64'b0010010111000101101000101001011100100110000001101010010111011101; end
            14'd6040 : begin out <= 64'b1010010011100000001010001100011110101000101000101010100000011000; end
            14'd6041 : begin out <= 64'b1010100010110100000110000110000000101010011011001001010010001010; end
            14'd6042 : begin out <= 64'b0010010111000000000111010110001000100011111010111010101110000001; end
            14'd6043 : begin out <= 64'b1010100001010000001010001110011010100100001011001010100101001110; end
            14'd6044 : begin out <= 64'b0010101010001011000101100011001100100111010100000010101111001110; end
            14'd6045 : begin out <= 64'b1010001001100110101010111001001010101000111101010010101110010000; end
            14'd6046 : begin out <= 64'b1010000101111110101001100010100100101000111110010010100000000000; end
            14'd6047 : begin out <= 64'b0010000011100100001010111011101000100101010100001010100010010100; end
            14'd6048 : begin out <= 64'b1010101110011010001010000001111100101010110101111001010011001100; end
            14'd6049 : begin out <= 64'b1010000010100101001001110001010010100111010101000010011001001101; end
            14'd6050 : begin out <= 64'b1010101101110001101001110110111100101000101110111010101100000101; end
            14'd6051 : begin out <= 64'b1001110000010011000010101010111100101001111001101010001101001101; end
            14'd6052 : begin out <= 64'b1010101001000000101010010011010010101001010111100001110001000100; end
            14'd6053 : begin out <= 64'b1010000101010011001001110100001010100010110111101010011111111100; end
            14'd6054 : begin out <= 64'b0010000101000101101010000010010100101010011011011010101000101111; end
            14'd6055 : begin out <= 64'b1010000101100010001001001011010100100010001001000010001100000001; end
            14'd6056 : begin out <= 64'b0010101000011010101010111100111110101000110111010001110111010000; end
            14'd6057 : begin out <= 64'b0010100111011111001000101010101100100010011010010001111101110011; end
            14'd6058 : begin out <= 64'b0010100101100001001010111010000110101010010111110010010010100110; end
            14'd6059 : begin out <= 64'b1010101100111111101010111111100110101010101110110010011000110001; end
            14'd6060 : begin out <= 64'b1010100010000101101010100101111000101000010111010010101011101100; end
            14'd6061 : begin out <= 64'b0010011110111011101001110110111010101010101000100010001010010111; end
            14'd6062 : begin out <= 64'b0010011011011011001010101010010110101000101000101001111001111011; end
            14'd6063 : begin out <= 64'b1010101001110001101010011101011110101000010001110001111001101101; end
            14'd6064 : begin out <= 64'b1010101111010110101010000001110100101011001000010010011010000110; end
            14'd6065 : begin out <= 64'b0010101111101110001001011010001000100110111100001010100011111101; end
            14'd6066 : begin out <= 64'b1010101010111010101010101011000000101100010011010010100001001111; end
            14'd6067 : begin out <= 64'b0010101101011111001010101100110100101010010011110010100001100010; end
            14'd6068 : begin out <= 64'b0010101110110110001010000110000010101010100101000010010110110100; end
            14'd6069 : begin out <= 64'b0010101000011101001010001100100110101010110011011010001000010001; end
            14'd6070 : begin out <= 64'b0010011100001101001010010000111110100000010100001010101101111110; end
            14'd6071 : begin out <= 64'b1010010000000001001010011111010010101010011010101010010101111011; end
            14'd6072 : begin out <= 64'b0010011000101111101001001000000010100111011111000010011010111000; end
            14'd6073 : begin out <= 64'b0010100001100001001001001001011100100010011101001001111110001110; end
            14'd6074 : begin out <= 64'b0010001101110001101010001111001000101010101100011010000101111101; end
            14'd6075 : begin out <= 64'b0001010110001010001010000011000010011101101111010010101011011010; end
            14'd6076 : begin out <= 64'b0010000110100000101010110101001110100101011100110010100110010110; end
            14'd6077 : begin out <= 64'b1010010010011010101001000111101100100110110110011010001100010100; end
            14'd6078 : begin out <= 64'b0000111000101010101000010100110010100101110110001001110000011101; end
            14'd6079 : begin out <= 64'b1010100000100100101000001111010010100111100011011010100110011101; end
            14'd6080 : begin out <= 64'b1010011100011000001010001111000010101010111000101010101111010110; end
            14'd6081 : begin out <= 64'b0010001101101111001010100010010100100000001001000001111100100000; end
            14'd6082 : begin out <= 64'b1010101000011010000111101011100110011011111100000010100000110010; end
            14'd6083 : begin out <= 64'b0010011111110111101010011111111000101000100101110010010011001101; end
            14'd6084 : begin out <= 64'b1010101100001000101010011011101010011101110011111010100101110100; end
            14'd6085 : begin out <= 64'b0010001101000011101010111110000010101001100001111010101010101100; end
            14'd6086 : begin out <= 64'b1010101101110010001010000101010110011010110000111010011100111001; end
            14'd6087 : begin out <= 64'b1010100111000010001010101110001000101000100000010010100100011111; end
            14'd6088 : begin out <= 64'b0010100100010101001010011100100000101010110100010010101011001010; end
            14'd6089 : begin out <= 64'b1010001000000011101001101110011100101000010010110010000000110101; end
            14'd6090 : begin out <= 64'b0010001100100101001010110011010110100110111110100010100100001100; end
            14'd6091 : begin out <= 64'b0010101111000111001010100110110000101000011000111010101111000110; end
            14'd6092 : begin out <= 64'b1010101110001110101010101100101110011011010100101010011111000110; end
            14'd6093 : begin out <= 64'b1010100010111000101001111100100110101001100110111010011110110101; end
            14'd6094 : begin out <= 64'b0010101000111100101010111000100000101010101100001010010100100001; end
            14'd6095 : begin out <= 64'b1010100000001111001010110111111000101010111110100010011010110101; end
            14'd6096 : begin out <= 64'b1010101001000101001010111110001010101010100110110010000110001011; end
            14'd6097 : begin out <= 64'b1010101111110110001010110011110100100110101011101010100111011101; end
            14'd6098 : begin out <= 64'b0010100011111100001010010010100100100110000011101010101110010011; end
            14'd6099 : begin out <= 64'b0010100101110101101000110000000000101000001110010010011001011101; end
            14'd6100 : begin out <= 64'b1010100111000100101010000110000110100100001101101010100110010011; end
            14'd6101 : begin out <= 64'b0010110000000000001010010111001000101001111111010010100000011100; end
            14'd6102 : begin out <= 64'b0010011111111100101010000001001100101010010011111010000001000110; end
            14'd6103 : begin out <= 64'b0010010111010000000111101100101010101001111010001001111111101010; end
            14'd6104 : begin out <= 64'b1001111010110000101001000001010100101000101111011010010010011010; end
            14'd6105 : begin out <= 64'b0010101000100110001001010010000010101010110011001001110000001011; end
            14'd6106 : begin out <= 64'b1010100100101110101001011011000100100010011010000010010100101110; end
            14'd6107 : begin out <= 64'b1010011100011001001001110111100110101011011100000010100001110010; end
            14'd6108 : begin out <= 64'b1010011011110101001010011000101000100100110010001010010111010111; end
            14'd6109 : begin out <= 64'b1010101011000101001000010010010000100101100110101010100001000111; end
            14'd6110 : begin out <= 64'b1001111000001101101001111010011010101001010000101010100011000111; end
            14'd6111 : begin out <= 64'b1001110101010100101001011000100010100101101001100010100111001010; end
            14'd6112 : begin out <= 64'b1010000011010111101000000101000100100011010000110010010111000101; end
            14'd6113 : begin out <= 64'b1001110101011110001010100001010100100111111010000010010001101011; end
            14'd6114 : begin out <= 64'b0010100101010110001010011100111010101010110111100010001101010101; end
            14'd6115 : begin out <= 64'b0001110101111101101010101011010100101000010110111010100011110111; end
            14'd6116 : begin out <= 64'b0010001100100011101000110000001000100101000100001010101110111000; end
            14'd6117 : begin out <= 64'b1010010000100011101010010111010110100111011101001010101001011000; end
            14'd6118 : begin out <= 64'b0010101001010011101001011011101110100111000001100010100010001001; end
            14'd6119 : begin out <= 64'b1010100000001001001010101001110000101011001010110010010000100010; end
            14'd6120 : begin out <= 64'b0010000011000110001010011110010010101010001001110010001110110101; end
            14'd6121 : begin out <= 64'b0010100110100101001001100111010000100011100100001010100000111000; end
            14'd6122 : begin out <= 64'b1010100010100101101010001000111000101010000011011001001000010011; end
            14'd6123 : begin out <= 64'b0010101010010111101001110101100010100111100111111001111100011011; end
            14'd6124 : begin out <= 64'b1010010000101010101001110000100000100101001101101010010011010101; end
            14'd6125 : begin out <= 64'b1010001001000010001010001001111010100110110011100010101001111001; end
            14'd6126 : begin out <= 64'b1010011110101110001001111111001000011010110111011010101011110011; end
            14'd6127 : begin out <= 64'b1010100111110011001010101110110100101000100100011010110000001001; end
            14'd6128 : begin out <= 64'b0010010001111011001010010001011010010011100010000010100100111101; end
            14'd6129 : begin out <= 64'b0010100011001011101010001100101010100100111000100010100111010000; end
            14'd6130 : begin out <= 64'b1010101100100111001010110111000100101000011001011010010011001110; end
            14'd6131 : begin out <= 64'b1010101000100111000111100101000110011101001111011010010010101011; end
            14'd6132 : begin out <= 64'b0010011000000100000110100001010110101010001010110010001111100110; end
            14'd6133 : begin out <= 64'b1010100110101010101001000111010100001111100101010010010000010001; end
            14'd6134 : begin out <= 64'b1010100111100011001010100111011110100111111001011010011011010110; end
            14'd6135 : begin out <= 64'b0010100110101001101001110001100100101010100110000010010000010110; end
            14'd6136 : begin out <= 64'b0001011001011110001010111010100000100111000111101010101011000101; end
            14'd6137 : begin out <= 64'b0010100001100000001001010010011110000101111101000010100110101000; end
            14'd6138 : begin out <= 64'b1010010111100010001000000011110100101001000101111010011100000101; end
            14'd6139 : begin out <= 64'b0010011111101100001001111000100010101000000000100010100011001111; end
            14'd6140 : begin out <= 64'b0010100001110001001000110111100100100010000111001010100000001011; end
            14'd6141 : begin out <= 64'b0010000000101011001010101101010000100100101000000010011010001010; end
            14'd6142 : begin out <= 64'b0010101000010111000100000100100110011100100001100010001100001011; end
            14'd6143 : begin out <= 64'b0001100000000111101001011011100110100100101011010010010111011010; end
            14'd6144 : begin out <= 64'b1001111110010000101010100101100100100101011010111010011011111101; end
            14'd6145 : begin out <= 64'b1010010100000100101010110011110100101011001110001010011001101111; end
            14'd6146 : begin out <= 64'b0001011110011100001010110011101000100100011010001001110111000101; end
            14'd6147 : begin out <= 64'b1010101010100001000111000010110000100111011010111010100100110000; end
            14'd6148 : begin out <= 64'b0010100001000000101010101010100000011101100100111010101110111100; end
            14'd6149 : begin out <= 64'b1010101111010110001010001110000010101001000010100010101000001111; end
            14'd6150 : begin out <= 64'b0010100101011111101001101111010110100011001000001010010001111100; end
            14'd6151 : begin out <= 64'b1010100010110001101001011000011010100011101000110010100001010001; end
            14'd6152 : begin out <= 64'b0010000101011011101010010101001000101011101000100010100010110011; end
            14'd6153 : begin out <= 64'b0010100111101010100110101000010100101000000100011010101001111100; end
            14'd6154 : begin out <= 64'b0010010110110101101001011001101000100011000101100010100001011000; end
            14'd6155 : begin out <= 64'b1010101010101101101001111001110010100010001100110010100110011010; end
            14'd6156 : begin out <= 64'b1010110000011001001010010011111100101001110011010010101110001101; end
            14'd6157 : begin out <= 64'b0010011110010011101001011011101100101010101101100010010110111001; end
            14'd6158 : begin out <= 64'b0010100010100111001011000100001100101000011000100010100111111101; end
            14'd6159 : begin out <= 64'b1010101000000011101010101101111110101000010111100010101001001000; end
            14'd6160 : begin out <= 64'b1010001111101101101010111100101000100111001101110010000011010001; end
            14'd6161 : begin out <= 64'b0010100010001101001010010110100100101001101001100010101110110011; end
            14'd6162 : begin out <= 64'b0010100000100000101010000111010100100101100011101010110000000110; end
            14'd6163 : begin out <= 64'b1010101001100001001010110101010010101010110000100010010101000101; end
            14'd6164 : begin out <= 64'b1010100110000010101001111000101000101000110111000010010000110010; end
            14'd6165 : begin out <= 64'b0010010000010000101001000100001000101010001110110010100100100110; end
            14'd6166 : begin out <= 64'b0010100111010010101000000001000110101001011001010010100110100100; end
            14'd6167 : begin out <= 64'b0010011101011010001001000110101110101001010010101010100011000001; end
            14'd6168 : begin out <= 64'b1010000111110101101010110101110100100011011101100010100010010001; end
            14'd6169 : begin out <= 64'b1000111110011011101010010010000110100110100111101010010110011011; end
            14'd6170 : begin out <= 64'b1010011001110010101000110011001010100110111101110010010101111001; end
            14'd6171 : begin out <= 64'b0010011110101110101001011001101000010100010001100010101010011111; end
            14'd6172 : begin out <= 64'b0001100010010100001010111110000110101000001011111010100001000000; end
            14'd6173 : begin out <= 64'b1001101011111100101011000100001010100011100011000010100001111111; end
            14'd6174 : begin out <= 64'b1010100111101100001001100110000000100010101110011010101101010001; end
            14'd6175 : begin out <= 64'b0010100111011110001001111101100010011011111111101001100011100100; end
            14'd6176 : begin out <= 64'b1010101001101010001001110110100010101001110000101010100001110101; end
            14'd6177 : begin out <= 64'b1010011011111101001000001110001100011000100010110010101010101101; end
            14'd6178 : begin out <= 64'b1001111001101010001010011111101100101000110100011010100110101111; end
            14'd6179 : begin out <= 64'b0010100001110111001011000001001010101001110111000010010000100000; end
            14'd6180 : begin out <= 64'b0010100010011101101001000011011110100100011100011010010010011101; end
            14'd6181 : begin out <= 64'b1010011101000101101001001000001110101010110001111010100100100111; end
            14'd6182 : begin out <= 64'b0010011001101111001010011011101100101011111110110010101110111111; end
            14'd6183 : begin out <= 64'b0001110101010000001000011001100110101001101110110001010011100101; end
            14'd6184 : begin out <= 64'b0010010100011101001010100100110100101001100011111010101011000101; end
            14'd6185 : begin out <= 64'b1010101111100111001001101011101100101000000111100010100001111110; end
            14'd6186 : begin out <= 64'b0001110111101101001000100111110100101010011001010010010111001110; end
            14'd6187 : begin out <= 64'b0010101100110011000111101111111010100101011101100001100100000101; end
            14'd6188 : begin out <= 64'b1010100010001111001010010010001100100110110111011001101010101000; end
            14'd6189 : begin out <= 64'b0010010101011100101001010111100010101010001000010010000101011111; end
            14'd6190 : begin out <= 64'b0010101110011001001001001101010100100101111011110010101110000011; end
            14'd6191 : begin out <= 64'b0010000100001110001000110010011000101000001110101010100000011100; end
            14'd6192 : begin out <= 64'b1010100011001000001010101010110110101011011101011001000001110111; end
            14'd6193 : begin out <= 64'b0010100010101001101010110101100100100110010110100010100110110000; end
            14'd6194 : begin out <= 64'b0010100001011110001010111100010010101001110000100010000001100010; end
            14'd6195 : begin out <= 64'b1010110000110100000111001010011100100101110110111010011111100101; end
            14'd6196 : begin out <= 64'b0010100111111111001000110001011010101011011011001010110000000000; end
            14'd6197 : begin out <= 64'b1010100100001100101001001000110100101000111011111001110010001110; end
            14'd6198 : begin out <= 64'b1010010001101000001010100000001110101011001101101010010111011001; end
            14'd6199 : begin out <= 64'b0010010011010111101010101100011110101010100011011010100100111111; end
            14'd6200 : begin out <= 64'b0010001111101010101000011110011110011111111010111010101010011000; end
            14'd6201 : begin out <= 64'b1010100111101111001010000110000110101010001001100010010000101111; end
            14'd6202 : begin out <= 64'b0010010110100011101010111111010010010000011111100010010010101110; end
            14'd6203 : begin out <= 64'b1010101110111101001001101101110100100110101000010010010010100101; end
            14'd6204 : begin out <= 64'b1010100011010000001010010111101110101010000111101010000011011100; end
            14'd6205 : begin out <= 64'b1010011000101111001010101000110010100000101100001010011010010111; end
            14'd6206 : begin out <= 64'b0010101001100001101010110001111010100101100101000010101101010011; end
            14'd6207 : begin out <= 64'b1010101001101000100100001100010100101001011101010010100001101010; end
            14'd6208 : begin out <= 64'b0010001011000111101010101110110110101010000010010010101101100101; end
            14'd6209 : begin out <= 64'b0010101010111100101001001010101010101000111011111010100110111010; end
            14'd6210 : begin out <= 64'b0010010010011001000111111110000100101010001000010001011011110011; end
            14'd6211 : begin out <= 64'b0010010111000010101001010101011000100110001101111010000000100001; end
            14'd6212 : begin out <= 64'b1010101010001001000011100101001110101000011100101010101010111001; end
            14'd6213 : begin out <= 64'b1010101000100110001010000100100000100110001101111010100100110010; end
            14'd6214 : begin out <= 64'b1010010001011100001010101101111110100000110001111010010010111010; end
            14'd6215 : begin out <= 64'b1010001001011001101000010110010100101010001001000010100111111100; end
            14'd6216 : begin out <= 64'b1010101011011100000111100010100000101000100100000001010110001100; end
            14'd6217 : begin out <= 64'b0010100101011000101001001001101110101100000100010010101011001011; end
            14'd6218 : begin out <= 64'b0010010001000000101011000101100010100101110011110010100010111101; end
            14'd6219 : begin out <= 64'b0010010000111010000111011011001100101010101110010010011101101001; end
            14'd6220 : begin out <= 64'b1010011011010000101010011101111100100110010001101010100101101110; end
            14'd6221 : begin out <= 64'b0010010000011010001001011011011000100111000011101010100100101111; end
            14'd6222 : begin out <= 64'b1010101100101001001001100010001100100000010100001010011011110000; end
            14'd6223 : begin out <= 64'b1010000011110110101010101100101100101011011011110001111111000001; end
            14'd6224 : begin out <= 64'b0010011000000100001010010110011110100110110110100010101001110000; end
            14'd6225 : begin out <= 64'b0010101101100000101001100111010010101010000110100001101111011111; end
            14'd6226 : begin out <= 64'b0010011011000100000111111010111000100000001001110010011011101001; end
            14'd6227 : begin out <= 64'b0010010111100000001001000011011100011101101001000010100010010101; end
            14'd6228 : begin out <= 64'b1010011001010101101001011111010010101010111100101010010011000010; end
            14'd6229 : begin out <= 64'b1010010010000011001010011100110100100100010010101010100001101011; end
            14'd6230 : begin out <= 64'b0010010000001111000010010001111010100110001011010010100001010010; end
            14'd6231 : begin out <= 64'b0010010110010000101001100110100000100101110110011001011110100011; end
            14'd6232 : begin out <= 64'b1010011100011000000111110011100000101001111100110001111101110100; end
            14'd6233 : begin out <= 64'b0010101101001001001010111000011110101001111111010010100100110011; end
            14'd6234 : begin out <= 64'b0010101100001010101010110101000000011101111011011010101110001111; end
            14'd6235 : begin out <= 64'b1010010111011000001001011011110100101010011110000010010111110001; end
            14'd6236 : begin out <= 64'b0010101010101101001011000111000010100010000000111010101011111011; end
            14'd6237 : begin out <= 64'b0010100010111100001000111100010010101011000110110010100010011000; end
            14'd6238 : begin out <= 64'b1010010010110010100110010110101010101000100100010010000001000101; end
            14'd6239 : begin out <= 64'b0010101000010110101001001000000000101000011001001010010101010110; end
            14'd6240 : begin out <= 64'b1010011001011000101001000100100110100100100100100010001111000101; end
            14'd6241 : begin out <= 64'b0010100011011000001010001001111110101010100101111010101000010111; end
            14'd6242 : begin out <= 64'b1010100111100100101001001110111000011011111001111010100101011101; end
            14'd6243 : begin out <= 64'b1010101011110100001010011010111110101000000001100010010001000111; end
            14'd6244 : begin out <= 64'b1010010100110110101010100110100010101000010011001010100010101111; end
            14'd6245 : begin out <= 64'b1010100010100000001010110010110110101000000100011010011000001111; end
            14'd6246 : begin out <= 64'b0010100000011101001010001111101010100100000110100010100011000011; end
            14'd6247 : begin out <= 64'b1010011100111011001000101101011100101011101100101010100001100100; end
            14'd6248 : begin out <= 64'b0010001101111011001001111100010010100000011110010001111100110000; end
            14'd6249 : begin out <= 64'b0010110000011111001010000100110010101001000001010001110111111000; end
            14'd6250 : begin out <= 64'b1010101000110000101010011110111100100001010111110001100110110001; end
            14'd6251 : begin out <= 64'b1010100110010101001010110010001010101000011111101010011110011110; end
            14'd6252 : begin out <= 64'b0010100001011110001000001011110110011100010011110010100000101010; end
            14'd6253 : begin out <= 64'b1010100100011111100101001110000010101011101011101010001100111101; end
            14'd6254 : begin out <= 64'b1010101001000111001010100110101110100111011100001010101010101111; end
            14'd6255 : begin out <= 64'b1010001011101010001001010001010100101001001111100010101000111111; end
            14'd6256 : begin out <= 64'b0010011101101110101001110100100010100001101001101010011100001111; end
            14'd6257 : begin out <= 64'b1010100000000101101001110101001000101001100010010001111010000011; end
            14'd6258 : begin out <= 64'b1001101101101011101010101110100100100111111110101010100111001001; end
            14'd6259 : begin out <= 64'b0001110011100100001010110001010110101000100000111010010101101001; end
            14'd6260 : begin out <= 64'b0010101000010000001010100000111000101001100001001010010100111100; end
            14'd6261 : begin out <= 64'b0000110010111101101000001100010110100101011010110010010110101101; end
            14'd6262 : begin out <= 64'b0010100110100100101001011010000110101011001010001010010000001001; end
            14'd6263 : begin out <= 64'b0010011111101111101001011110100000101010101100110010011011101111; end
            14'd6264 : begin out <= 64'b1001111101010000001001111000011100101010101100000010100010100010; end
            14'd6265 : begin out <= 64'b1010000101100010001010001011011010101010100011111010101101100100; end
            14'd6266 : begin out <= 64'b1010010011101010001001110111010100100101001110001010011011000101; end
            14'd6267 : begin out <= 64'b0010000101000011001010110011100010011111011110011010010111100110; end
            14'd6268 : begin out <= 64'b0010101001011101101010111101011100100100001100001010010001011010; end
            14'd6269 : begin out <= 64'b1010010101101010001010110001000110101010100111010010010000110101; end
            14'd6270 : begin out <= 64'b0010001110011100101001101001001000101000010110100010100111111010; end
            14'd6271 : begin out <= 64'b1010101010111000101010010101000010011100111101000001011111101001; end
            14'd6272 : begin out <= 64'b0010011100000100001010101101110010101000100101000010100011010001; end
            14'd6273 : begin out <= 64'b0010011010000111101001101000001000100110111101011010100110101110; end
            14'd6274 : begin out <= 64'b1010010011010000001000011000111110101010101110111001110101011001; end
            14'd6275 : begin out <= 64'b1001011111011100001010111101000000101011100110001010101011000101; end
            14'd6276 : begin out <= 64'b0010001101110011101001000100100110101000001100110010010111100100; end
            14'd6277 : begin out <= 64'b0010101000101000001000111110011000100110011000001010100010100100; end
            14'd6278 : begin out <= 64'b1001100100111101101000111111111000100011011010111010101101010101; end
            14'd6279 : begin out <= 64'b1010010011101001001010000010110110101001000001100010100010011011; end
            14'd6280 : begin out <= 64'b0010101010101100001001001000010010010111100000011010010110010000; end
            14'd6281 : begin out <= 64'b0010001110000100001010110010110010101011000110000010101101011011; end
            14'd6282 : begin out <= 64'b1010100011011111001000100110110010101000010111101010010000110001; end
            14'd6283 : begin out <= 64'b1010101101111011101010010111101010100010110010111010100101110001; end
            14'd6284 : begin out <= 64'b0010011110100011101010010010101010101011101101000010001010010110; end
            14'd6285 : begin out <= 64'b1010100000110100001001100111001010101000001110000010001101010101; end
            14'd6286 : begin out <= 64'b0010011000011001101000110010110110001111010000111010100101110010; end
            14'd6287 : begin out <= 64'b1001111111101101101010110011101110101000000100000010100101110100; end
            14'd6288 : begin out <= 64'b0010101010001010000101010101111100100111110000100010001110101110; end
            14'd6289 : begin out <= 64'b0010011110101001001010001101101110101010100001100010101011101110; end
            14'd6290 : begin out <= 64'b1010001111110111101001110100000100101011000100100010101101001010; end
            14'd6291 : begin out <= 64'b1010010111101010001001000011111110100100000001110010010101010101; end
            14'd6292 : begin out <= 64'b0010010001111101101010001111101100101000111000100010101111011010; end
            14'd6293 : begin out <= 64'b0010011101100100001001010110000100100111000000110010101011111011; end
            14'd6294 : begin out <= 64'b0010010101100111101001100110000100101010111100111010101101000101; end
            14'd6295 : begin out <= 64'b0010000110111100001010111000110000101001000111101010101101101101; end
            14'd6296 : begin out <= 64'b1010100000000100001001110101001110101000100110110010100111010001; end
            14'd6297 : begin out <= 64'b0010101011000100101000110010111100101000101000100010010000000000; end
            14'd6298 : begin out <= 64'b0001110010110011101010110000111000101010100000011010100010110010; end
            14'd6299 : begin out <= 64'b0010100101111001101010111100111110011110111110101001101010110000; end
            14'd6300 : begin out <= 64'b0010100110010011100110101001100100010100101011011010101100101001; end
            14'd6301 : begin out <= 64'b1010100001110011001000001000011100011110110110101010101000100100; end
            14'd6302 : begin out <= 64'b0010010111011010001001001001101010101001100110100010101111000100; end
            14'd6303 : begin out <= 64'b0010101011001011101000100110100100100001001011011010000000001110; end
            14'd6304 : begin out <= 64'b0010100101100110100111100001010100101010101100101010101011011010; end
            14'd6305 : begin out <= 64'b1010100110110000001000011100100110100100011101100010101001110110; end
            14'd6306 : begin out <= 64'b1010010001000110101010010100011000100111111110101010100000110011; end
            14'd6307 : begin out <= 64'b1010101111000101001010000000110000100101100010001010001100101111; end
            14'd6308 : begin out <= 64'b0010101010011000101001101011100010101000011111101010001100010101; end
            14'd6309 : begin out <= 64'b0010100100000101101010001010011010101011101010000010000001111100; end
            14'd6310 : begin out <= 64'b0001010000110010001010100101110110101000010111000001110000001100; end
            14'd6311 : begin out <= 64'b1001110111010101101000001001000010101001100000100010101001010101; end
            14'd6312 : begin out <= 64'b0010001011110011101011000001011110101011000100011010100001101001; end
            14'd6313 : begin out <= 64'b1010101100001011001000100011111110101000110010101010010100010100; end
            14'd6314 : begin out <= 64'b1010101100111000001000000011101010101010110110011010101110010110; end
            14'd6315 : begin out <= 64'b1010000000101001001010101101100010101000111010011010101000001101; end
            14'd6316 : begin out <= 64'b0010011111001010000100010110001100100000001000001010000111000000; end
            14'd6317 : begin out <= 64'b1010101010001100001010101001000010100001100011100010011000000011; end
            14'd6318 : begin out <= 64'b0010110000111011001010111011111110011011110110111010101010010110; end
            14'd6319 : begin out <= 64'b1010011100110110001001100111101000100111010001001001110100000101; end
            14'd6320 : begin out <= 64'b0010101110101011101010101110101110100011110101111010101100011110; end
            14'd6321 : begin out <= 64'b0010100010100001001001100101111010101001010111011010100010011110; end
            14'd6322 : begin out <= 64'b1010010101101001001010101011110100100101010000000010011111001111; end
            14'd6323 : begin out <= 64'b1010101101000100101010011100000000011110011111000010000001011000; end
            14'd6324 : begin out <= 64'b1010100101111101101001111111001110101000000000010010101001101101; end
            14'd6325 : begin out <= 64'b1010010010111101101001100001111100101010011110101001101000010011; end
            14'd6326 : begin out <= 64'b1001111100000100001010000000110100101000100011111010010011010010; end
            14'd6327 : begin out <= 64'b1001010101000110001001011000011110100100110101011010100101011011; end
            14'd6328 : begin out <= 64'b1001011100101011100111110010001110100001101111100010010111111111; end
            14'd6329 : begin out <= 64'b1010001110011001001001101100110100100101001001011010101111100101; end
            14'd6330 : begin out <= 64'b0010100111010101001000001110001110100111010011110010000100111101; end
            14'd6331 : begin out <= 64'b0001101101011010100111101010100110101001111001011010101010001101; end
            14'd6332 : begin out <= 64'b1010100101111000001000010000110110101011100011100010100110010101; end
            14'd6333 : begin out <= 64'b1010101101010110000111010110010110101010000100110010100010010000; end
            14'd6334 : begin out <= 64'b1010100010101110101010111001110010101001111001100010100111010101; end
            14'd6335 : begin out <= 64'b0010011001001010100111001011000010101011110011101010101101000101; end
            14'd6336 : begin out <= 64'b1010010011111000001010000100101110101001011111010010100110011001; end
            14'd6337 : begin out <= 64'b0010101100111001001010101001100010100011001100111010000100010010; end
            14'd6338 : begin out <= 64'b0010100111111110101000100011100100100001011101111010010010100000; end
            14'd6339 : begin out <= 64'b0010011011110101100110110100111110101010100001101010100000101010; end
            14'd6340 : begin out <= 64'b1010010001001000101010011010100010100100110101110010100010100111; end
            14'd6341 : begin out <= 64'b1010100010101011001010011001011000100101010011001010100001100110; end
            14'd6342 : begin out <= 64'b1001111100111001001001000000101000100110000111100010100110101001; end
            14'd6343 : begin out <= 64'b1010101000100101100110101011000110101010011001101010011110000000; end
            14'd6344 : begin out <= 64'b1010010011001011101001110000011110101011001010001010100010111101; end
            14'd6345 : begin out <= 64'b1010101001111111101001100001111010100100100100010010100100011101; end
            14'd6346 : begin out <= 64'b0010100000001001001010101000110110101001011111000010100101010010; end
            14'd6347 : begin out <= 64'b1010100111010010001010111100100100101010111101110001111010111101; end
            14'd6348 : begin out <= 64'b1010101101011001001000011111000110101000001000001010100110001110; end
            14'd6349 : begin out <= 64'b0010101100100100001001011101000000100001111011101001110000000011; end
            14'd6350 : begin out <= 64'b1010101010100100100111000010010100101000001100011010101110011001; end
            14'd6351 : begin out <= 64'b1010101000110011001000101010001110100001011001001010100011010000; end
            14'd6352 : begin out <= 64'b1010101101011100101001000101010100100011010011000010100010101110; end
            14'd6353 : begin out <= 64'b1001010100001010001010101011010000011100001101100010011100101000; end
            14'd6354 : begin out <= 64'b1010100110111000001010110000011000101010011100010010100001110000; end
            14'd6355 : begin out <= 64'b0010101101000100001001100011011000100000111101101010011000111001; end
            14'd6356 : begin out <= 64'b0010101111101000101010010100110010100110111010000010100000010011; end
            14'd6357 : begin out <= 64'b0010100001111001101000100010100110101010000011001010100011110100; end
            14'd6358 : begin out <= 64'b1001101101110011101010100101100010101010000001010010100000000010; end
            14'd6359 : begin out <= 64'b0010001111000001100111001111001100101010000111110010101100000000; end
            14'd6360 : begin out <= 64'b1010100001011010100111010100010110100100001110110010101001111101; end
            14'd6361 : begin out <= 64'b0010011100111010000101110011100000101100010100011010010001110110; end
            14'd6362 : begin out <= 64'b1010100001010010001000101101100010100101001000111010100110100110; end
            14'd6363 : begin out <= 64'b0010101010000110001010100000101100101000010111010010101111001100; end
            14'd6364 : begin out <= 64'b1010011001111110000111011011010010101010001111111010101110001101; end
            14'd6365 : begin out <= 64'b1010101100000101101000101001100010100010000000111010100101011001; end
            14'd6366 : begin out <= 64'b0010101111001100101010001110110000100010100100111010010000010000; end
            14'd6367 : begin out <= 64'b0010100110011011001001000000100000101000100110101010000001010111; end
            14'd6368 : begin out <= 64'b0010011101010001001010100011101000101001000111011010100011010100; end
            14'd6369 : begin out <= 64'b0001110100101101101010010000111010100111111100110010000001101110; end
            14'd6370 : begin out <= 64'b0010100001100001101010011000100110100001000110011010011010001110; end
            14'd6371 : begin out <= 64'b1010000011001010101010001100101110100011010001101010010001111110; end
            14'd6372 : begin out <= 64'b1010100000000111101001011110011000101010101101010001111110101001; end
            14'd6373 : begin out <= 64'b1010101110100011101010101101100010101001101010000010011110110000; end
            14'd6374 : begin out <= 64'b1010010111011111001010101101110010101010010111000010101011101101; end
            14'd6375 : begin out <= 64'b0001100110101110001001101101100010100100111101110010100111001011; end
            14'd6376 : begin out <= 64'b0001110000010001101010001001000010011101111101110010101000100100; end
            14'd6377 : begin out <= 64'b1010010101100110000100111011000000011110011011000010011011000011; end
            14'd6378 : begin out <= 64'b0001011000110001001000011000101110101011011101000010001011110101; end
            14'd6379 : begin out <= 64'b1010100111000011100101011110101110101001001110111010011000100001; end
            14'd6380 : begin out <= 64'b0010001111100111001010001101110110100100100001010010100110110010; end
            14'd6381 : begin out <= 64'b0010100101111110001001010110000000100101111110101010100001110100; end
            14'd6382 : begin out <= 64'b1010100011101101001010110111001000101001100001111010010100111110; end
            14'd6383 : begin out <= 64'b1010010010001011001001101110000010101001011011110010100010111100; end
            14'd6384 : begin out <= 64'b0001111010101100101000001000001100101001101000100010100000100111; end
            14'd6385 : begin out <= 64'b0010011110000000001010000111000110100101000001100010011110010110; end
            14'd6386 : begin out <= 64'b0010001101110010001001001101010010010101101100111010101010100011; end
            14'd6387 : begin out <= 64'b1010010110100111001000011100011010100110101010100001010011101101; end
            14'd6388 : begin out <= 64'b0010000000000110001010101110111010101001111011101010000111111100; end
            14'd6389 : begin out <= 64'b0010010010100001001010010101100110100110110011000010101100010011; end
            14'd6390 : begin out <= 64'b1010001011111011101010010110011100101011110011011010101000110011; end
            14'd6391 : begin out <= 64'b0001100100001001101000000011000110101010011110011010100110000011; end
            14'd6392 : begin out <= 64'b1010101010011110000111111101010110100100110000000010100000101000; end
            14'd6393 : begin out <= 64'b0010100011110000001010111010011100011110111100000010101100100101; end
            14'd6394 : begin out <= 64'b1010011001100111001010101011010100101011100110000010011001110101; end
            14'd6395 : begin out <= 64'b0010001100100101101010111110010100100010001110111010010100100010; end
            14'd6396 : begin out <= 64'b0010001111100110001000011110001110101001100001001010100010110101; end
            14'd6397 : begin out <= 64'b0010100111011001101001100000011010100101000000110001001000110100; end
            14'd6398 : begin out <= 64'b0010100110100011001001110111100010100110010111011010010110000111; end
            14'd6399 : begin out <= 64'b0010100000110001001000110001011000101000011010001010010001010000; end
            14'd6400 : begin out <= 64'b0010100011001111001010101011101010101011001101101010000011001011; end
            14'd6401 : begin out <= 64'b0010100100000101001010000111010110011110111100111010101001001110; end
            14'd6402 : begin out <= 64'b1010001011001100001010101011000000011100001010101001010111111011; end
            14'd6403 : begin out <= 64'b1010010101111011001010111011101000101010100100000010101001100101; end
            14'd6404 : begin out <= 64'b0010010100110011000100000110000110010110001111011010100010010001; end
            14'd6405 : begin out <= 64'b0010010000000101001010110010100010010100101010000010100100100010; end
            14'd6406 : begin out <= 64'b1010011111101110001001010001101010101010000101111010000110100110; end
            14'd6407 : begin out <= 64'b0010101101111001100100010010000010011000000011011010101100011000; end
            14'd6408 : begin out <= 64'b0010011100001100000111011101011010010000101001011010101110010101; end
            14'd6409 : begin out <= 64'b0010100001100010000011101100001100101000100000111010101010100000; end
            14'd6410 : begin out <= 64'b1010001100010111001010011110101100100110001011110010010011001110; end
            14'd6411 : begin out <= 64'b1010100011110100101010100011000010100111010011101010011100111000; end
            14'd6412 : begin out <= 64'b1010001000111100101010010110111010101011111111001010101101100100; end
            14'd6413 : begin out <= 64'b1010101010111011101001000111010110101011000011010010001010110001; end
            14'd6414 : begin out <= 64'b0010011000010011101010110011100000101010000010111010001111001000; end
            14'd6415 : begin out <= 64'b0001111110011000101010111100110000101100000000111010010010111110; end
            14'd6416 : begin out <= 64'b0001110011101001101010010111110010101001000100101010100011100100; end
            14'd6417 : begin out <= 64'b1010011011000011001001011000000010100001000001010010011001100001; end
            14'd6418 : begin out <= 64'b0010010101001110101001010010100010101001001001011010100110001101; end
            14'd6419 : begin out <= 64'b1010010110111011101010011001000010101001010001001001100101101101; end
            14'd6420 : begin out <= 64'b0010100001111010001010010111110000100110011100010010101000100010; end
            14'd6421 : begin out <= 64'b0010100111100111001001110001100010100110101011001010101110011111; end
            14'd6422 : begin out <= 64'b0010101010000000001001101111011000100111111011000010101001101110; end
            14'd6423 : begin out <= 64'b0010101010100101001001000011001000101100000001001001101100001111; end
            14'd6424 : begin out <= 64'b0010010100100010001010011111100000100111100101110010100100100001; end
            14'd6425 : begin out <= 64'b0010001111010100101010000100011010100010011110111010011100001000; end
            14'd6426 : begin out <= 64'b1010011000110111001010010010010010101011001000101010100100100110; end
            14'd6427 : begin out <= 64'b0010100001001110101010011001111110101010100110100010101101010011; end
            14'd6428 : begin out <= 64'b1010100110100101101000000010001100100011011000011010000100011001; end
            14'd6429 : begin out <= 64'b0010001110111000001001100001000100100010111011101010101100010101; end
            14'd6430 : begin out <= 64'b0010100010001100001010100011100010101001110101110010001000011101; end
            14'd6431 : begin out <= 64'b1010101110010110001010100101001110101010011101000010010011000000; end
            14'd6432 : begin out <= 64'b0010000000001110101000011111011100100111010111100010101010001111; end
            14'd6433 : begin out <= 64'b0010101110010000101010100101010100100100010111111010101111111100; end
            14'd6434 : begin out <= 64'b0010011001110111100111001011011100101001101111011010010001111101; end
            14'd6435 : begin out <= 64'b1010100011111101101001101001100100101011100010101001101010100111; end
            14'd6436 : begin out <= 64'b1010101000110100001001000101110010101000000110000010101011001010; end
            14'd6437 : begin out <= 64'b1010100000001100001010000110110000100001111011100010011100101011; end
            14'd6438 : begin out <= 64'b0010100111111110001010111111011000011011000100110001111000010111; end
            14'd6439 : begin out <= 64'b0010001100001010000111110111101000101001010111011010101110011111; end
            14'd6440 : begin out <= 64'b0010010101101111101010000101100100101001000001110010100110001101; end
            14'd6441 : begin out <= 64'b0001010000010011001000101011111110011001011101001010100010001000; end
            14'd6442 : begin out <= 64'b1010000001000011001001011110000110100010101000000010101011101101; end
            14'd6443 : begin out <= 64'b0010000111100010001000000001011100101011111100000001111111101001; end
            14'd6444 : begin out <= 64'b0010101100100010001001001110101000100100101001110010001110111001; end
            14'd6445 : begin out <= 64'b1010010001110010001001101100101110101001010100100010101111100010; end
            14'd6446 : begin out <= 64'b1010101000001011000111101101010010101011011011011010000100010111; end
            14'd6447 : begin out <= 64'b1010101101111010101001010001011100101011010011101010010101011110; end
            14'd6448 : begin out <= 64'b1010010101111011001001110110010000101000010111000001111100010111; end
            14'd6449 : begin out <= 64'b0010101000001001001010000100111110100110111000111010011001010010; end
            14'd6450 : begin out <= 64'b0010101011011111101010000101010010101011100111110010100001001110; end
            14'd6451 : begin out <= 64'b0010101110101110001001100001100110100101011010011010010000010001; end
            14'd6452 : begin out <= 64'b0010010100101100001001101001001110101011110110100010101000010111; end
            14'd6453 : begin out <= 64'b1010100100110000101001010101110110100011101110111010101000100111; end
            14'd6454 : begin out <= 64'b1010010000011011000111100101010100101010000000011010100101000010; end
            14'd6455 : begin out <= 64'b0010010001001010101010011111101000101011110001101010101000100011; end
            14'd6456 : begin out <= 64'b1010011111010101101010001000110010101000011100011010101011111100; end
            14'd6457 : begin out <= 64'b0010101000100001101000010101011100100101101110001010010111111110; end
            14'd6458 : begin out <= 64'b1010000110100101001001111001100100010110110000111010011100100101; end
            14'd6459 : begin out <= 64'b1010100110101010101010110101001010101011110101011010101010111111; end
            14'd6460 : begin out <= 64'b0001100010011010000110010111110010101011111000101000000110111111; end
            14'd6461 : begin out <= 64'b1010000010000000001010000111001010101010001011100010001011100101; end
            14'd6462 : begin out <= 64'b1010100000000110001001110101011110100100001110001010000010010000; end
            14'd6463 : begin out <= 64'b1010100101010001000111111111111100101010001001111010101110111000; end
            14'd6464 : begin out <= 64'b1010100101111001101000110111011100101000000110011010101000100110; end
            14'd6465 : begin out <= 64'b0010100110101100001010001100101100101011010011101010101011100001; end
            14'd6466 : begin out <= 64'b1010100111101111001010111111110010100111000000011010000100111110; end
            14'd6467 : begin out <= 64'b1010011001101110101010011011010100100111001111100010101111011011; end
            14'd6468 : begin out <= 64'b0001100011100010101010111110010110100100010111000001110001101000; end
            14'd6469 : begin out <= 64'b1010010011001100001010011000000010101000100010001010101001101010; end
            14'd6470 : begin out <= 64'b1010010101101001000111110110011000101010111110000001100101110010; end
            14'd6471 : begin out <= 64'b1010011111100010001010011011011010101011100000111010000000011111; end
            14'd6472 : begin out <= 64'b1010100000001000101001011001011100101001101011100010100111011110; end
            14'd6473 : begin out <= 64'b0010101010001001001001100011110110101000000111100010100100110001; end
            14'd6474 : begin out <= 64'b0010100000000111001001000101111010100110110010010001110101001101; end
            14'd6475 : begin out <= 64'b0010101011011101001010111010011110101010001111001010100110010000; end
            14'd6476 : begin out <= 64'b1010101100100011001001001001000110010110111111010010101111111001; end
            14'd6477 : begin out <= 64'b0010010101101100001010111001111010101011100011000010010011101100; end
            14'd6478 : begin out <= 64'b1010100010000011100111111111011110101010111011101010101010101000; end
            14'd6479 : begin out <= 64'b0010101101111011001010110010010110100010110111110001110100010100; end
            14'd6480 : begin out <= 64'b0010000000011101001010100001010010011111010010001010000010000010; end
            14'd6481 : begin out <= 64'b0010010000000001001001000100000000100001011010111010011110111100; end
            14'd6482 : begin out <= 64'b0010101101111100101010110011101000000000110111111001110011000100; end
            14'd6483 : begin out <= 64'b1010100000011101001010100101110100100100111010011010001111100100; end
            14'd6484 : begin out <= 64'b1010101010001011101010101101110110011110011001001010100000001011; end
            14'd6485 : begin out <= 64'b0010011101100101101010100110000100101010111001101010100001111111; end
            14'd6486 : begin out <= 64'b1010100011100100001001011101101100101011011110011010100110111011; end
            14'd6487 : begin out <= 64'b0010011010110100101010010111100010011101111000011010010111001110; end
            14'd6488 : begin out <= 64'b0010010010000000001001001010100100100010100110010010010100101100; end
            14'd6489 : begin out <= 64'b1010011001011100001010011010111110011111110100000010101010000101; end
            14'd6490 : begin out <= 64'b1010000111111000000111101011001000101000010111010010100001010110; end
            14'd6491 : begin out <= 64'b1010100010110101101000011000001110100110100101111010011001110001; end
            14'd6492 : begin out <= 64'b0010011101111110001000101011000010101010001111001001101010100000; end
            14'd6493 : begin out <= 64'b0010100011001000101010111001111110011000111100001010010001010100; end
            14'd6494 : begin out <= 64'b1010100110000100101011000000101110101001011101101010101100110110; end
            14'd6495 : begin out <= 64'b1010001010011001001010000011100000100100011011111010100001101110; end
            14'd6496 : begin out <= 64'b0010011001110111101010100000000000100101001110101010011100110110; end
            14'd6497 : begin out <= 64'b1010010010001111101010110000100110101001001100100010010100001000; end
            14'd6498 : begin out <= 64'b1010011001001101100110110000100010101010001001100010001110111100; end
            14'd6499 : begin out <= 64'b0010101001101110101010001000101100010100100010000010100100000101; end
            14'd6500 : begin out <= 64'b0010101110010101101010000010111110010100000101110010101011011001; end
            14'd6501 : begin out <= 64'b1010011110110000001010101000001110100001011000000010010101001100; end
            14'd6502 : begin out <= 64'b1010100100011110101010001111010100100100100111111010100000011111; end
            14'd6503 : begin out <= 64'b0010101010101000101010000100101000100111000111110010100000100011; end
            14'd6504 : begin out <= 64'b1001101111100001101001101000010000100100110001001010011010011010; end
            14'd6505 : begin out <= 64'b0010101101101110001001100110111010011111111000000010101000100110; end
            14'd6506 : begin out <= 64'b0010100101000101001010101001101100101011111000000010101111000001; end
            14'd6507 : begin out <= 64'b0010101011011011101010000001110110101000000111100010100111111011; end
            14'd6508 : begin out <= 64'b0010101000101100001001010010110000101001101011001010101110001111; end
            14'd6509 : begin out <= 64'b1010000000111101001010000010010100101010100000111010011110010001; end
            14'd6510 : begin out <= 64'b0010011110111010101010110011011100100101000001111010010100001011; end
            14'd6511 : begin out <= 64'b0010010001110100001010010011110000101001011100011010010011001111; end
            14'd6512 : begin out <= 64'b0010010111000110001010011111000000100100011111001001110100011111; end
            14'd6513 : begin out <= 64'b1010101111001111001001011001100100100101110001101010011010010111; end
            14'd6514 : begin out <= 64'b1010101111100101001010010011111100100101101000101010010010001110; end
            14'd6515 : begin out <= 64'b0010100010001010001010010111001100101000000000001010001000011001; end
            14'd6516 : begin out <= 64'b0010010110010110101010010011110000101000000001101010001001111010; end
            14'd6517 : begin out <= 64'b0001100100111100101010010000100010101010000100111010011111000111; end
            14'd6518 : begin out <= 64'b0010100011101111101010001111101100100111010111000010101001000100; end
            14'd6519 : begin out <= 64'b0010001010011011001010000011011000101001110111011010011101101100; end
            14'd6520 : begin out <= 64'b0001111101000011101010110001110100101010110000100010100110100101; end
            14'd6521 : begin out <= 64'b1010000111000100100101101111001000101011100010000010011000101000; end
            14'd6522 : begin out <= 64'b0010101110111100001010000101110010010111001001100010001110000010; end
            14'd6523 : begin out <= 64'b0010011111011100001001001010001100101011010001100001101101010001; end
            14'd6524 : begin out <= 64'b0010101111111110001001100010101000101000101110000010011110111101; end
            14'd6525 : begin out <= 64'b1001111101011011001000100100010000001100100100110010100111110010; end
            14'd6526 : begin out <= 64'b0010010001000101001001100100100100100110001000000010000111010011; end
            14'd6527 : begin out <= 64'b0010101111100101001010100010111010101000011111110010101010111111; end
            14'd6528 : begin out <= 64'b1010100010110101101001000101100100101000111110101010101101001011; end
            14'd6529 : begin out <= 64'b0010001011101100001010010101000100100100100001111010011100111100; end
            14'd6530 : begin out <= 64'b1010100111101110001010101101011100011010011000101001111111101001; end
            14'd6531 : begin out <= 64'b0010011011001100101010010011100110101010011110111010011000101011; end
            14'd6532 : begin out <= 64'b0010100110110001101010000101111110100011101100101010100111000110; end
            14'd6533 : begin out <= 64'b1010101100110000100011110111110100101010111100111010101010000010; end
            14'd6534 : begin out <= 64'b1010001010000111101000010001100010011000101001111010011010011010; end
            14'd6535 : begin out <= 64'b0010011010100101100101100001011100101001110111000010001000010110; end
            14'd6536 : begin out <= 64'b0010100011010001001001101010010010101000110110111010010111100010; end
            14'd6537 : begin out <= 64'b0010100000111101001001011101111000101011011010110010101110100100; end
            14'd6538 : begin out <= 64'b1010100110111110100101100010111100011111001000110010100110000100; end
            14'd6539 : begin out <= 64'b1010100011110011001001011101110000100010111100011010101111101111; end
            14'd6540 : begin out <= 64'b1010100100110000001010110000010000010001000111010010101001111110; end
            14'd6541 : begin out <= 64'b0010010010101000101010101011111110101000111000010010001010110000; end
            14'd6542 : begin out <= 64'b0001110100110111101010101100010100001001111111011010100110001111; end
            14'd6543 : begin out <= 64'b1010010101010011101010000100010000100101100110001010010110111111; end
            14'd6544 : begin out <= 64'b0001110000100111001000110001110000101000010010111010000110001011; end
            14'd6545 : begin out <= 64'b0010100111010000101010000101110110100110000001010010000001011001; end
            14'd6546 : begin out <= 64'b1010001011110011101010001011010100101010100111111010100011100001; end
            14'd6547 : begin out <= 64'b1010101100110110001001010000111000100110111000000010001100010100; end
            14'd6548 : begin out <= 64'b0010011111000101001010010001110010100100000001000001101101000000; end
            14'd6549 : begin out <= 64'b1010101001101100001010000010110010100100011000011010000011011101; end
            14'd6550 : begin out <= 64'b1010101100010011100111101110101110100011111110000010100010101111; end
            14'd6551 : begin out <= 64'b0010010110100100000110000001000110100111000010111010001101110000; end
            14'd6552 : begin out <= 64'b1010101001001010101010011110110110101000111100001010000101111011; end
            14'd6553 : begin out <= 64'b1010100011000001101010000100001100100110100111010010101011111011; end
            14'd6554 : begin out <= 64'b0010101101001001001010100101110010011100010000011010101100100101; end
            14'd6555 : begin out <= 64'b1010101110101100001010001000110110100011101111111010101011111110; end
            14'd6556 : begin out <= 64'b1010000110010011101000000011100110101010111101011010100101100010; end
            14'd6557 : begin out <= 64'b1010011001000010001010101011100110100000000000100010100110110100; end
            14'd6558 : begin out <= 64'b0010101010100101101001011000100010101011110100011010010100110110; end
            14'd6559 : begin out <= 64'b0010100010100100101010101010111110100110110101000010101000010111; end
            14'd6560 : begin out <= 64'b1010100000111110001010011001010100101100000010100010011111000100; end
            14'd6561 : begin out <= 64'b0010100011101110101001100011100100100010001110011010011010111001; end
            14'd6562 : begin out <= 64'b0010010001000100100111001011010000101010100101001010100000110110; end
            14'd6563 : begin out <= 64'b1010010101101001101010000110000010101011000101111010101011101110; end
            14'd6564 : begin out <= 64'b1010001100000101101010000000011010100111111111011010100110000100; end
            14'd6565 : begin out <= 64'b0010001111100010101010101001001100101010010100000010100000010001; end
            14'd6566 : begin out <= 64'b1010101011001110001010011100011010100110010110101010101000000101; end
            14'd6567 : begin out <= 64'b1001110011110000101010011111011000100010010111001010010100011100; end
            14'd6568 : begin out <= 64'b0001110100010111001010000000010110101000101100010010101110111100; end
            14'd6569 : begin out <= 64'b1010101110101101101000101110110000100101000001000010000011110010; end
            14'd6570 : begin out <= 64'b0010100011001000100101110001011000101001100001000010100111111111; end
            14'd6571 : begin out <= 64'b0010011101001101001010011011101010101000101101010010101000111000; end
            14'd6572 : begin out <= 64'b0010011101000001001010010100111000101000101000011010010000110001; end
            14'd6573 : begin out <= 64'b1001110000001101101010011001000000101010010101010010101100100011; end
            14'd6574 : begin out <= 64'b0001011100100001101010110011100110010100000000101001111100101010; end
            14'd6575 : begin out <= 64'b0010010111111111101010011111010110100110111010001010100110101111; end
            14'd6576 : begin out <= 64'b0010011110110101101001110110000010101010100001001010100010110000; end
            14'd6577 : begin out <= 64'b1010001001101000101001011111111000100001101001101010101011110000; end
            14'd6578 : begin out <= 64'b1001110011101100001010111011100110100101001111101001111111000101; end
            14'd6579 : begin out <= 64'b0010100111100100100101001100011100101011101110111010100011010010; end
            14'd6580 : begin out <= 64'b1010011011011100001001001011001110100000000011111010010110100001; end
            14'd6581 : begin out <= 64'b1001000110101001101001101110010000101010110111001010010110110001; end
            14'd6582 : begin out <= 64'b1010011101000010001010111011110110101010100011001010100101111001; end
            14'd6583 : begin out <= 64'b0010010101010101000111000010010000011000010100001001111010111011; end
            14'd6584 : begin out <= 64'b1010001110001111101010111101110010100110111101101010010101111011; end
            14'd6585 : begin out <= 64'b0010101011011000101010001100010110100110011111110010010010101010; end
            14'd6586 : begin out <= 64'b0001010111000011101010110010001010101001111110001010010100110110; end
            14'd6587 : begin out <= 64'b1010101011010001101010011011110100101001110111011010011100001110; end
            14'd6588 : begin out <= 64'b0010010100000101001001101100000010100100100110011001001011110111; end
            14'd6589 : begin out <= 64'b1010001010000110001000111010101110100110010110110010101000110001; end
            14'd6590 : begin out <= 64'b1010101111001001101001001000001000011100101111110010101011001000; end
            14'd6591 : begin out <= 64'b1010010010110011101000010011000110100110001011111010101111100011; end
            14'd6592 : begin out <= 64'b1010100010011110001001001111010010101001110101110010101100000010; end
            14'd6593 : begin out <= 64'b1010101100011001001001110100001000100101010011101010100011100001; end
            14'd6594 : begin out <= 64'b1010101100110011101010001000010110101000110111111010100101000010; end
            14'd6595 : begin out <= 64'b1010100011001000001001010001000000101000100000010010001110010001; end
            14'd6596 : begin out <= 64'b1010101100100110001010111100001100101000101101101010101100001011; end
            14'd6597 : begin out <= 64'b1010101000010101001001001010010110100001001101111010010100111001; end
            14'd6598 : begin out <= 64'b0010100101001011101010110010110100100111000100000010010101110100; end
            14'd6599 : begin out <= 64'b1010001010111000000110101101110010001101000001101001010010011000; end
            14'd6600 : begin out <= 64'b0010101001001110001010111111001010101010111011100010100000010010; end
            14'd6601 : begin out <= 64'b1010100110101010001001110010010100011110110111000010010110100010; end
            14'd6602 : begin out <= 64'b1001110011011010101010000101110100100110010011111001101100101111; end
            14'd6603 : begin out <= 64'b1010101000010110101001000011111110101011000000010010010000000111; end
            14'd6604 : begin out <= 64'b0010100110000011101000001011000100100111010101110010011111111011; end
            14'd6605 : begin out <= 64'b0010010011110000001010000010110000100100001001101010100000111100; end
            14'd6606 : begin out <= 64'b1010100111001000101001010010010100100111101001001010100111010011; end
            14'd6607 : begin out <= 64'b0010100100101110101010001001011010100001011000111000110101110100; end
            14'd6608 : begin out <= 64'b0010000100101011100100111011001010100000101011001010011100110000; end
            14'd6609 : begin out <= 64'b1010101011110110101001111001110000101011011000100010100010111001; end
            14'd6610 : begin out <= 64'b1010011101001011001001101110001100100101010111110010100111110110; end
            14'd6611 : begin out <= 64'b1010000101001000101000000011111000101000110101111010100011010000; end
            14'd6612 : begin out <= 64'b0010101001101010001001001011000110100011111011000010010110001010; end
            14'd6613 : begin out <= 64'b0010101101011111101001101100000010101000110001101010000100101101; end
            14'd6614 : begin out <= 64'b0010010010111000101010010000111100101011011101100010001111101011; end
            14'd6615 : begin out <= 64'b1010010111000001000111011010010110010100001101010010100010101101; end
            14'd6616 : begin out <= 64'b1010100010001111001000011001010010101001111110111010101000111101; end
            14'd6617 : begin out <= 64'b1010000000011011101010101110011110101000111000111010100101110011; end
            14'd6618 : begin out <= 64'b1010101101111011101010010111011110100010001001011010000111110101; end
            14'd6619 : begin out <= 64'b1010010001110101001000110000010000010011110001110010001001101000; end
            14'd6620 : begin out <= 64'b0010010101110100101010000110011000101010101101001010101110101010; end
            14'd6621 : begin out <= 64'b1001110000100010101010001000100000100111000000100010011101100100; end
            14'd6622 : begin out <= 64'b0010001111110010001010000001001100101011110011110010101111010011; end
            14'd6623 : begin out <= 64'b0001110101110100001010001001110000101001000001110010100111001101; end
            14'd6624 : begin out <= 64'b0010100110011000001001110101110010100010111011000010011101110000; end
            14'd6625 : begin out <= 64'b1001011101001110001010001101000010010001000111101010011111011001; end
            14'd6626 : begin out <= 64'b0010101100101010001010011101010000011110001010110010101100110001; end
            14'd6627 : begin out <= 64'b1010100010000101101010010001110000100100100111000010010110101000; end
            14'd6628 : begin out <= 64'b1010010011101011001010010000101100100111100000000010100010101101; end
            14'd6629 : begin out <= 64'b1010011111101111001010111010101010101011010000011010100010101110; end
            14'd6630 : begin out <= 64'b0010010110001111001010010011110000100110010100110010100111111000; end
            14'd6631 : begin out <= 64'b1010010111100011101001110100100010101001000011010010100010100101; end
            14'd6632 : begin out <= 64'b1001101001101001101010011001000000101011000101000010100110101011; end
            14'd6633 : begin out <= 64'b1010101101001000001010111000110100101010110001010010011111010001; end
            14'd6634 : begin out <= 64'b0010011110000110101000001111110110011100110011000010011001110100; end
            14'd6635 : begin out <= 64'b1010011010100011101010000001000000101011001100100010011111010001; end
            14'd6636 : begin out <= 64'b0010100110010110101010011110001110100001001010001010011010001100; end
            14'd6637 : begin out <= 64'b0010101011110111001001000001000110101001101000100010000110001110; end
            14'd6638 : begin out <= 64'b0001111001100101101000011010111110011101001011100001111111000011; end
            14'd6639 : begin out <= 64'b1001111001101001000111101101011100101000001101010010101110110100; end
            14'd6640 : begin out <= 64'b1010100101011101100011101100010010011011010001000010100010110000; end
            14'd6641 : begin out <= 64'b0010100111110110001000010010000100101000000100010010000001110000; end
            14'd6642 : begin out <= 64'b0010011111101001001010000101100100101000100100111001000111001101; end
            14'd6643 : begin out <= 64'b1010011110001100101010100100000110100100000001100010001001010111; end
            14'd6644 : begin out <= 64'b0010000110110110001010010101111000100110000010000010100100110100; end
            14'd6645 : begin out <= 64'b0010101110101011101001111000001000100101111110011010001000100001; end
            14'd6646 : begin out <= 64'b0010010001111101001010011011111100100101001101001010100001010001; end
            14'd6647 : begin out <= 64'b1010010100011011000111000000110000011100000100101010000110000111; end
            14'd6648 : begin out <= 64'b1010100111000100101010110011111010100110100111000010101011001010; end
            14'd6649 : begin out <= 64'b0001100101011110000110000110001000101011010101000010100011111011; end
            14'd6650 : begin out <= 64'b1010011011111010101001110001000110101000101000011010010101000010; end
            14'd6651 : begin out <= 64'b0010101010011101101010011011011100011110111110000010100101001011; end
            14'd6652 : begin out <= 64'b1000100001001110001001111110010100100001000111001010101001001001; end
            14'd6653 : begin out <= 64'b0010101100010011001010010111111100100101000011110010100101010110; end
            14'd6654 : begin out <= 64'b0010011111101010001000011001010000101010011110010001110111110011; end
            14'd6655 : begin out <= 64'b1010001010011100101010101001110110101000001011000010100110000011; end
            14'd6656 : begin out <= 64'b1010101010101101101001100110110010011110011001100010100110001111; end
            14'd6657 : begin out <= 64'b1001100001001100001010110000111110101000010011000010101110011110; end
            14'd6658 : begin out <= 64'b1001010100011110101000011101010100100011101001111010100110111000; end
            14'd6659 : begin out <= 64'b1010100100000110001010111111111010101011000010100001100010111000; end
            14'd6660 : begin out <= 64'b1010000111111010101010010011001110101000000110011010101110011000; end
            14'd6661 : begin out <= 64'b1010101000110011001001011101010100101010110111110010101010111111; end
            14'd6662 : begin out <= 64'b0010101011101101101000011011011110101001101010101010010010010110; end
            14'd6663 : begin out <= 64'b1010101010011101001001001100110110100011001111110010101100111001; end
            14'd6664 : begin out <= 64'b0010011000100101101001010101101100101010111000100010011011111010; end
            14'd6665 : begin out <= 64'b0010010101111101001001110110101110100110100000000010000110110011; end
            14'd6666 : begin out <= 64'b1010100001101001101001100001010010100110110101110010101010000010; end
            14'd6667 : begin out <= 64'b1010101100001101001010100011110000100100000110000010010001001111; end
            14'd6668 : begin out <= 64'b0010001000100011001001111110101110101001110100010010011010100010; end
            14'd6669 : begin out <= 64'b0010101000101100001001001110110100101011111100001010101101010001; end
            14'd6670 : begin out <= 64'b0010010101100001101001010000100000101000101111000010101100011000; end
            14'd6671 : begin out <= 64'b0010100010110110101001100011010100101010011101011010010000100110; end
            14'd6672 : begin out <= 64'b0010011010001011101001010101111110100111101100110010100000111011; end
            14'd6673 : begin out <= 64'b0010100110001100101010001101011110100101100110101001101010101011; end
            14'd6674 : begin out <= 64'b0010100011101010101001111111101110101010111011000010101111000010; end
            14'd6675 : begin out <= 64'b1010101100011101001010010110010100101001001000101010011001100011; end
            14'd6676 : begin out <= 64'b1010101001000010101010110001101000100011000010011010100111010110; end
            14'd6677 : begin out <= 64'b1010001100001010001010010111100010101001101101000010101111011011; end
            14'd6678 : begin out <= 64'b0010101011000011101010001101000000011000011100100010010000110011; end
            14'd6679 : begin out <= 64'b1010011101111101101001101000011110100000110001001010100100011111; end
            14'd6680 : begin out <= 64'b0001100110111110101010111110101110100101110111110010010100111110; end
            14'd6681 : begin out <= 64'b1010001100000111101001100101011010011101110010100010100101100010; end
            14'd6682 : begin out <= 64'b0001110100010111101001111110110000101000110001100001111010011101; end
            14'd6683 : begin out <= 64'b0001100001001001001010110000000000011001100000001010011010110010; end
            14'd6684 : begin out <= 64'b0010011011100000101010010111000110101010101001101010101011001000; end
            14'd6685 : begin out <= 64'b1010011010010011000110001110001000101000111110010010011111010100; end
            14'd6686 : begin out <= 64'b0010100110001110001010001111010100101000001011110010100000110001; end
            14'd6687 : begin out <= 64'b1010101001100110101010000111000010101011101001011010011100110100; end
            14'd6688 : begin out <= 64'b1010101110001010101010001100111110101011101100110010011101111001; end
            14'd6689 : begin out <= 64'b1010101111001110001001000001100000101011111010100010001000100111; end
            14'd6690 : begin out <= 64'b1001001110111100101001010010111000101011100111111010101000000100; end
            14'd6691 : begin out <= 64'b1010100010001001101000100100101110100010010101011010001111010011; end
            14'd6692 : begin out <= 64'b1010101100100011101010111100111000100010101000000010010110110001; end
            14'd6693 : begin out <= 64'b1010100100000110100111111111110010100110011010100001100110110110; end
            14'd6694 : begin out <= 64'b0010100010110010001010001000001100101011001111001010010011111001; end
            14'd6695 : begin out <= 64'b1010101000111000101010010010000010101011000001110010000110100001; end
            14'd6696 : begin out <= 64'b1001100000000001101010001101111110100100001011000010010110111100; end
            14'd6697 : begin out <= 64'b0010101011111101100100000010010010100110110000100010011010111010; end
            14'd6698 : begin out <= 64'b1010001100111100101000100111010110100101101001010001110001011001; end
            14'd6699 : begin out <= 64'b0010011101110001101010010000110000100110001011010001111110100110; end
            14'd6700 : begin out <= 64'b1010001001000101101001000011010000101001100110101010100110011111; end
            14'd6701 : begin out <= 64'b1010101001010000101010010101101110100100101001011010101101011000; end
            14'd6702 : begin out <= 64'b1010100101000001101001101101110110100101100111110010010110100010; end
            14'd6703 : begin out <= 64'b0010101011011010001010100111110100100101011111101010011011010101; end
            14'd6704 : begin out <= 64'b0010000100100101101010111110101010101000001100000010100110110011; end
            14'd6705 : begin out <= 64'b0010100000011000100111000000100000101001111011000010100110101011; end
            14'd6706 : begin out <= 64'b1010100100111101001010010100001100101000001100111010011001111101; end
            14'd6707 : begin out <= 64'b1010101100010011101000110100001100101001001100111010110000010000; end
            14'd6708 : begin out <= 64'b1010010110011001101010011111101100101011101001110010001000011001; end
            14'd6709 : begin out <= 64'b1010100010000001101010111011000110101011100100000010100110000101; end
            14'd6710 : begin out <= 64'b0010101110001100101010110000000100100101001000000010101001000000; end
            14'd6711 : begin out <= 64'b0010100110010001101001000110010000100011100001100001010101010000; end
            14'd6712 : begin out <= 64'b1010101110010110100111110110011100101001100001000010101111011111; end
            14'd6713 : begin out <= 64'b1001101111111100001010111101100000011010011100101010000101100100; end
            14'd6714 : begin out <= 64'b0010101100001100101001111110010100100001111101110010010010000111; end
            14'd6715 : begin out <= 64'b0010001000100000100110100001000100100000110100111010000100010101; end
            14'd6716 : begin out <= 64'b0010011010110110101010111110111010101001001100011010101100110110; end
            14'd6717 : begin out <= 64'b1010010011101000000101101110000110101000100011001010100101101100; end
            14'd6718 : begin out <= 64'b1010001011110111101010111000110100101010110100011010010100111100; end
            14'd6719 : begin out <= 64'b1010100100101010001010010101100000100111010100110010101000001100; end
            14'd6720 : begin out <= 64'b0010011100100001101010100001111100101001011011101010101100000110; end
            14'd6721 : begin out <= 64'b0010011101010101001001000101101010100110101101111010101101111010; end
            14'd6722 : begin out <= 64'b1010011110101110001010000011100110100111011010011010011100001100; end
            14'd6723 : begin out <= 64'b1010000011010101101010001110100110101011001111111010001101111001; end
            14'd6724 : begin out <= 64'b0010001000110100101001000101011110101011010111110010101100011111; end
            14'd6725 : begin out <= 64'b0010010000100110000111110110110110100010111001011010101101001011; end
            14'd6726 : begin out <= 64'b1010010100111100101001110001101010101010001110100001011011111000; end
            14'd6727 : begin out <= 64'b0010101011101001001010010111000000010110111101111010100001101100; end
            14'd6728 : begin out <= 64'b1010011011010111001010100101100000101000010101010010000100100011; end
            14'd6729 : begin out <= 64'b1010000110011111001000000111110100101010101101100010011100111001; end
            14'd6730 : begin out <= 64'b1010100110100100000100110111000100010110100000101010000100101001; end
            14'd6731 : begin out <= 64'b1010101101010101101000001011001000100101111011100010010101000111; end
            14'd6732 : begin out <= 64'b1010011101000110000111011001110010101001101110110001010011110010; end
            14'd6733 : begin out <= 64'b0001101111001001101010011011111110100111110111001010101110011101; end
            14'd6734 : begin out <= 64'b1010100001011111101010001000110010101011011011110010101110001110; end
            14'd6735 : begin out <= 64'b0001110010100011001010010111000100100111010000110010101000101110; end
            14'd6736 : begin out <= 64'b0010100001101111001010101001010110100100111011111010100110110100; end
            14'd6737 : begin out <= 64'b1010101010101011101010100100111010100101110100110010100110001101; end
            14'd6738 : begin out <= 64'b1010101001101110001000101111110000101001010000100010101011100010; end
            14'd6739 : begin out <= 64'b0010101011110110101010011001100010101100001010111010101111010000; end
            14'd6740 : begin out <= 64'b1010100011010111101010010100101100100100111100111010100101111001; end
            14'd6741 : begin out <= 64'b0010010001000001101010111011011110101001101101101001111111101011; end
            14'd6742 : begin out <= 64'b1010011000010101001001000111110110101010100000010010100000101110; end
            14'd6743 : begin out <= 64'b0000110001110111001000001000101110011101011011111010100010000011; end
            14'd6744 : begin out <= 64'b0010101110010100101010100001011010101001000110111010101101111001; end
            14'd6745 : begin out <= 64'b0010100100000010101001000011001000101000001010010010001011010110; end
            14'd6746 : begin out <= 64'b0001110001010100001001110010011010100011011010110010011011011110; end
            14'd6747 : begin out <= 64'b1010100011000111001010000110100010101010000010011010101110000101; end
            14'd6748 : begin out <= 64'b0010011111111010000111010110011110101001010001111001101101010010; end
            14'd6749 : begin out <= 64'b0010011011110101101010000011110110101010001110011010101100011110; end
            14'd6750 : begin out <= 64'b0010000011000110001010101001011010100111001101001010010000100010; end
            14'd6751 : begin out <= 64'b1010011100101101101010100101001010101001000111110010101011010000; end
            14'd6752 : begin out <= 64'b1001110010110001101010001101110000100110101001010010011000110001; end
            14'd6753 : begin out <= 64'b1010100010000000000110001001001100101010011001111001011110010001; end
            14'd6754 : begin out <= 64'b0010101011100100001010011111111100101001101110110010001111001000; end
            14'd6755 : begin out <= 64'b0010100110001111101010001011100010011100010100000001100101000010; end
            14'd6756 : begin out <= 64'b1010100001110111001001100011111100100010010101100010101011111111; end
            14'd6757 : begin out <= 64'b0010100010000110001010001011111110100010110110101001110100100100; end
            14'd6758 : begin out <= 64'b0010101001111010101001101001110000101011100001011010101011110100; end
            14'd6759 : begin out <= 64'b0001111111011101101010110001101000101010101111100010010101110010; end
            14'd6760 : begin out <= 64'b0001100010110110101001010000100010101000100001000010110000000101; end
            14'd6761 : begin out <= 64'b0010010100011010001000101011000010100110010010000010000000011010; end
            14'd6762 : begin out <= 64'b1010010110010011101001010001100100101011001001111010001001001101; end
            14'd6763 : begin out <= 64'b1010101010000010101010111001010110101000110011110010011100101000; end
            14'd6764 : begin out <= 64'b0010010001100101101010010010010100101000000111111010011011001100; end
            14'd6765 : begin out <= 64'b0001111101110010101010001000010000101011101010000010010001011010; end
            14'd6766 : begin out <= 64'b0010100000100100100110101000101010101010011100010010101001101010; end
            14'd6767 : begin out <= 64'b0010101100011000101010111100001010101000000110001010100110101001; end
            14'd6768 : begin out <= 64'b0010100101110100101010111011000100000000110010011010101011000000; end
            14'd6769 : begin out <= 64'b1010000000000010101000011001111110100001000110010010100100111001; end
            14'd6770 : begin out <= 64'b1010100011100010101010100001010110100101110101111010101000110110; end
            14'd6771 : begin out <= 64'b1010100111000001001010010111110100101010110111011001010000110110; end
            14'd6772 : begin out <= 64'b0010100110000001101000010111101110101011001010101010100010111100; end
            14'd6773 : begin out <= 64'b1010100111010010001010001011000110100111011111000010000000110111; end
            14'd6774 : begin out <= 64'b0010001010101011001001011111110010100011110011001010100010000000; end
            14'd6775 : begin out <= 64'b0010010001000010101010110011011110101001010000001001110000000001; end
            14'd6776 : begin out <= 64'b0010001101010011001001011011110100100011011111111001101010011111; end
            14'd6777 : begin out <= 64'b0010010101011010001010100111010110100010010001101010101110100001; end
            14'd6778 : begin out <= 64'b0010101010010111101001001010010000101010111111100010100111110000; end
            14'd6779 : begin out <= 64'b1010011010101100100110001111100110100000111001010001100001111010; end
            14'd6780 : begin out <= 64'b0010100001110001001000110000111110010111100001111010100000010111; end
            14'd6781 : begin out <= 64'b1010100101001101001001001010001110100001011101101010101010111100; end
            14'd6782 : begin out <= 64'b0001110001111010101010010001011000101001010110011010100000100100; end
            14'd6783 : begin out <= 64'b0010011100101110001000101001010010100010011000100010001101011101; end
            14'd6784 : begin out <= 64'b1010011000010001001010010101001000101011100100111010100110110001; end
            14'd6785 : begin out <= 64'b1010101010001110101001110101000110100100000110100010011001011000; end
            14'd6786 : begin out <= 64'b0010011011111010101010010100000010101000000110100010010110100101; end
            14'd6787 : begin out <= 64'b1010010101000110100110001110100000101010100000000010100000000100; end
            14'd6788 : begin out <= 64'b0010101101011011101001000011100010100101001111100010101100101001; end
            14'd6789 : begin out <= 64'b0010010100100111000111110111001100101000000011110010010010011110; end
            14'd6790 : begin out <= 64'b0010100111010010001001000100111110101010001110000010010100011100; end
            14'd6791 : begin out <= 64'b0010100000111001101010101001101110100011000101111010011110010001; end
            14'd6792 : begin out <= 64'b1010000010010110000111101111110110100110000111010010010111011111; end
            14'd6793 : begin out <= 64'b0010100010101101101001000111110000101100001101001001110011111011; end
            14'd6794 : begin out <= 64'b0001101111000011001000001011110000100111110101001010101011110111; end
            14'd6795 : begin out <= 64'b1010100010000100101010101111011110011110011000101010101000101010; end
            14'd6796 : begin out <= 64'b0010011000101111101010111101100110101011011010001010100011110101; end
            14'd6797 : begin out <= 64'b1010101011100101101010011101111100100110100010001010100110111111; end
            14'd6798 : begin out <= 64'b0010011111101001100111010111101100100010000011110010010101011001; end
            14'd6799 : begin out <= 64'b0010100000010011101001101001011110101000011111001010101111100101; end
            14'd6800 : begin out <= 64'b0010101010011111001010101011011000100100110000100010011101110010; end
            14'd6801 : begin out <= 64'b1010100111001001101010001111111000101001000110101010100101000111; end
            14'd6802 : begin out <= 64'b0010000101110111101001000110110010101000001111000010000000110101; end
            14'd6803 : begin out <= 64'b1010100000110110101000001110000100100001101111100010010001110001; end
            14'd6804 : begin out <= 64'b1001000000010011101010110001000100100101111011100010010001001101; end
            14'd6805 : begin out <= 64'b1010000100100111101001010001111110100110010011000010000111000011; end
            14'd6806 : begin out <= 64'b1010100101001000101010110000011000100111010010001010100110110100; end
            14'd6807 : begin out <= 64'b1010101011111111100111010101100100100010001000011010001000010101; end
            14'd6808 : begin out <= 64'b0001111010001011101010111001111010101001000111011010100101100110; end
            14'd6809 : begin out <= 64'b1001011110101110101010100111011010101001011011100010011011000001; end
            14'd6810 : begin out <= 64'b1001111000001110001001001011000100101010000000111000111110110110; end
            14'd6811 : begin out <= 64'b0001101110110000001001011010100010011101010100010010101010101011; end
            14'd6812 : begin out <= 64'b0010101100011010101001001111110010101000000100100010100110100010; end
            14'd6813 : begin out <= 64'b0010010111111000100111101101111010101010001111011010010011111010; end
            14'd6814 : begin out <= 64'b1010001010010111100100010101010000101000000011110010010010000100; end
            14'd6815 : begin out <= 64'b1010101011101001001010101110111110100101100100010001101001111011; end
            14'd6816 : begin out <= 64'b1010100001110001001010001000000110011100101000011001100111010111; end
            14'd6817 : begin out <= 64'b0001110101010010101010100001110000101000010010100010001100111001; end
            14'd6818 : begin out <= 64'b0010010011011111001010010100010010101010000100110001100110110111; end
            14'd6819 : begin out <= 64'b1010100111111000001010110000011110101010111010110010100010001110; end
            14'd6820 : begin out <= 64'b1010100101111011101010110001111100101001111100101010100001010101; end
            14'd6821 : begin out <= 64'b0010101001001000001010010000010100101001100100011010100001011000; end
            14'd6822 : begin out <= 64'b0001100000111111001010110101100110011100011110111010000111000111; end
            14'd6823 : begin out <= 64'b1010010111001000000110010011100110100111110000010010100010111100; end
            14'd6824 : begin out <= 64'b1010101111011110001010110101010000100110101001001010101000011101; end
            14'd6825 : begin out <= 64'b1010010001010011101001011010111010101011110100000010010101111111; end
            14'd6826 : begin out <= 64'b1010100011001000101001110101000110101000001101011010101010110110; end
            14'd6827 : begin out <= 64'b1010101000100011001010001010011100100110101100010010100111111010; end
            14'd6828 : begin out <= 64'b0010100000011011001001000001010110100111111100101010101001101001; end
            14'd6829 : begin out <= 64'b1010100000001100101010100000010110101011011010000001111110110001; end
            14'd6830 : begin out <= 64'b1010010111101100101001100000101100101011101101101010101011100000; end
            14'd6831 : begin out <= 64'b0010101000001011001010010111001010010001000000010010000100111010; end
            14'd6832 : begin out <= 64'b1010011000100111101010010011001100101001000100101010100001010011; end
            14'd6833 : begin out <= 64'b1010100100101011100100111111010110100000000000100010101100010010; end
            14'd6834 : begin out <= 64'b1010100111101111101001011011111110011111000011011010100100001100; end
            14'd6835 : begin out <= 64'b0000111100111111001010011000101100010011001111000010001110111010; end
            14'd6836 : begin out <= 64'b0010011001110001001001011101111010100000110001111010011010010001; end
            14'd6837 : begin out <= 64'b1010000001100001001001101110100010101010110000111010101100100110; end
            14'd6838 : begin out <= 64'b0010011100010000000101110110101100101001101000000010101111010001; end
            14'd6839 : begin out <= 64'b1010010000100110001001010000111000101001100000001010100100110000; end
            14'd6840 : begin out <= 64'b0010001001101100000011000001100110101001101011100010101111010001; end
            14'd6841 : begin out <= 64'b0010000001000010001010111001110100100101000010011010010001001010; end
            14'd6842 : begin out <= 64'b1010100001110100001010110010010000101001000100011010011111110101; end
            14'd6843 : begin out <= 64'b0010101110101011100111101111001100100000010000010010100010011101; end
            14'd6844 : begin out <= 64'b0010010101110001001010101011011100101010010010110010100000110011; end
            14'd6845 : begin out <= 64'b1010000100111100001010010111100100001111111110101001110001001101; end
            14'd6846 : begin out <= 64'b1010010001110100001001111010011000100111101101100010011101110001; end
            14'd6847 : begin out <= 64'b1010100111010100101010101011100000100110011010001010001100110111; end
            14'd6848 : begin out <= 64'b1010010000100100000111001010110110100101111001000010100000101110; end
            14'd6849 : begin out <= 64'b0010101001010100001001011110100110101001011010110010011110011110; end
            14'd6850 : begin out <= 64'b0010010111101100101010110100101010101011111110100010010010101001; end
            14'd6851 : begin out <= 64'b1010100000011000101010101101101100100101100101111010100011100001; end
            14'd6852 : begin out <= 64'b1010100000110101001000001010100000101011101101101010101001010010; end
            14'd6853 : begin out <= 64'b0010100101111000101000101001001010101010110110001010100001111000; end
            14'd6854 : begin out <= 64'b1010100010100110101001100001111110101011000011001010010011000011; end
            14'd6855 : begin out <= 64'b0010011001111101101010110111011000101010110000011010001100001001; end
            14'd6856 : begin out <= 64'b1010011001000100001001011101001110100110100110111010001011100011; end
            14'd6857 : begin out <= 64'b0010001001111010101000100010010110101000011001100010100110111001; end
            14'd6858 : begin out <= 64'b0001111010111101001001100111011010101011110111010001100111000001; end
            14'd6859 : begin out <= 64'b1010100000100001001010010101001000100010000001011010100000111000; end
            14'd6860 : begin out <= 64'b0010100000111001001001110110110100101001111011010010100101001001; end
            14'd6861 : begin out <= 64'b0010011011011011001000011111011110101000101000110010010011000011; end
            14'd6862 : begin out <= 64'b1010100110100010001010111010010010101001101101101010010110111101; end
            14'd6863 : begin out <= 64'b1010010110010001101000001110101010100010111101100010101011100011; end
            14'd6864 : begin out <= 64'b1010000001010111101001110110110000011111110001110001101001001001; end
            14'd6865 : begin out <= 64'b0010000111100010101001000111000010100111111000000010001010001011; end
            14'd6866 : begin out <= 64'b0010100101110011101001001110000100011001011110001010000110010001; end
            14'd6867 : begin out <= 64'b1010101101101001101010111100111110100101001010000010000101001011; end
            14'd6868 : begin out <= 64'b1010011000011111001010110001111010101010011000011010000111000100; end
            14'd6869 : begin out <= 64'b0010100011111011001010100100101010100110010111101010011100101001; end
            14'd6870 : begin out <= 64'b0010100011010100001010011001111000100000110111001010100111111010; end
            14'd6871 : begin out <= 64'b1010010010110110101000000000101100100001010011110010000100000011; end
            14'd6872 : begin out <= 64'b1010011000101010001010111000001110100000000101100010101001000101; end
            14'd6873 : begin out <= 64'b1010010111000001101010011111000000100100110000111010010010011010; end
            14'd6874 : begin out <= 64'b1010100000000101101010010000100100100111010110111001101001011111; end
            14'd6875 : begin out <= 64'b1010100001100110101010010111011100101001110001011010010101100110; end
            14'd6876 : begin out <= 64'b1010011100011011001000111000111010100000111000000010011100101000; end
            14'd6877 : begin out <= 64'b1010101111001000001000111101011110100001000110110010011111111110; end
            14'd6878 : begin out <= 64'b1001110100011010001010101100000110100111110111101010000111100110; end
            14'd6879 : begin out <= 64'b1010100111001110000100110000101110011000111111100010010001101111; end
            14'd6880 : begin out <= 64'b0010010110111001101000000000001000101001001010010010010011110100; end
            14'd6881 : begin out <= 64'b0010101001101101101001010110101100101000010110100010000001000010; end
            14'd6882 : begin out <= 64'b0010101110010000101000101111001110101001001110110010010001111000; end
            14'd6883 : begin out <= 64'b0010010100110100101010001001000000100001001101111010010100001101; end
            14'd6884 : begin out <= 64'b0010011100100011101010110101001010101011101010000010101100110010; end
            14'd6885 : begin out <= 64'b0010001010011101001010100010100110100110011000001001101100111010; end
            14'd6886 : begin out <= 64'b0010101000101100101010110111101100100111110010000010100000100100; end
            14'd6887 : begin out <= 64'b1010011000010111101011000000100010101001110101100001100010111110; end
            14'd6888 : begin out <= 64'b0001100010111011100111011001000010101011001111000010001111100100; end
            14'd6889 : begin out <= 64'b0010011101100101101000001001110110101010101111010010100000100111; end
            14'd6890 : begin out <= 64'b1010100100100110101010001101101000100000110100100010010001010001; end
            14'd6891 : begin out <= 64'b1010011101101110100111011110010100100111001101010010101011000011; end
            14'd6892 : begin out <= 64'b0010101011010101101010010100000000011111101000010010100000000010; end
            14'd6893 : begin out <= 64'b1010010010111111101010001000101010101000110101011010100101100001; end
            14'd6894 : begin out <= 64'b0010010000111011101010010100000110011100001101001010101101100101; end
            14'd6895 : begin out <= 64'b0010000010111001101000001100000000101011001110001001110100111010; end
            14'd6896 : begin out <= 64'b1010010001101110001000111101100010000001001000111010010111010010; end
            14'd6897 : begin out <= 64'b1010100100010001101011000000100010100100101101111010001101101000; end
            14'd6898 : begin out <= 64'b1010010101011110101001000111010100100111110100011010010110011001; end
            14'd6899 : begin out <= 64'b0010101001110011001010000011000000100111000111011010101011011001; end
            14'd6900 : begin out <= 64'b0001110110100101001000001111010100101010101010000001001111000010; end
            14'd6901 : begin out <= 64'b1010101100100000100111010101110010101010011001100010011011011111; end
            14'd6902 : begin out <= 64'b1010011001000111101010001100001100101010101101100010101010010001; end
            14'd6903 : begin out <= 64'b0010000111000111001001011010001100100111001101001010100000010011; end
            14'd6904 : begin out <= 64'b1010010011000111001010010100001010100100000100100010000011000010; end
            14'd6905 : begin out <= 64'b1010001111010001001000010110000100101001010001100001100000101010; end
            14'd6906 : begin out <= 64'b1001001100101110101000110011011110101001000010111010011111000111; end
            14'd6907 : begin out <= 64'b1010101101001111101000000110101110100011100100110010000000000000; end
            14'd6908 : begin out <= 64'b1001010111011111000110110000111110101010001010110010100000110010; end
            14'd6909 : begin out <= 64'b1010100011011001001001001110011010101000010111011010100000110010; end
            14'd6910 : begin out <= 64'b1001111001101010001000110001011110011111001011011010100111101100; end
            14'd6911 : begin out <= 64'b0010010011010000001000000110001010011100001011001010011010111111; end
            14'd6912 : begin out <= 64'b0010110000000001101010110011010010101011001001100010101101011111; end
            14'd6913 : begin out <= 64'b0010010101001001001010110010001010100110101000100010010011001100; end
            14'd6914 : begin out <= 64'b0010001011110011101010111100000100101000101001000010101100011101; end
            14'd6915 : begin out <= 64'b0010100100011011100101101000111100101000010110000010101101111111; end
            14'd6916 : begin out <= 64'b0001011110110101001001001010111000100000001011010010101000111000; end
            14'd6917 : begin out <= 64'b1010010010101000101010001110011010101001110111001010011011000000; end
            14'd6918 : begin out <= 64'b1010100011000110000110010100111110101001001100011010011010111111; end
            14'd6919 : begin out <= 64'b1010101110000010001001101100101000100010110001001010010000111010; end
            14'd6920 : begin out <= 64'b0010101010110001101010010101001110100111110011101010101000000000; end
            14'd6921 : begin out <= 64'b0010101011111000101010101010011100100111001100110010101110101001; end
            14'd6922 : begin out <= 64'b1010101111001000001010100000011100100101100100000010101101001011; end
            14'd6923 : begin out <= 64'b0010100000101011101001010100000110101011100001110001111111100100; end
            14'd6924 : begin out <= 64'b1010100111001110101000000011101010100101101010001010100000011101; end
            14'd6925 : begin out <= 64'b1010100011111100101010100001010110101011110000100010100111101101; end
            14'd6926 : begin out <= 64'b1010100010001110001001111111100010101010110010111010000010011110; end
            14'd6927 : begin out <= 64'b1010101011000111001001011110110010101011100001010010100111101111; end
            14'd6928 : begin out <= 64'b1010101110011001000110110101111010100110110100011001111000000111; end
            14'd6929 : begin out <= 64'b0010101000010110001010100110010000101000101100000010101101000111; end
            14'd6930 : begin out <= 64'b1010001001001100101010101111111100100111110000101010101010011100; end
            14'd6931 : begin out <= 64'b1010101110001110101010001111001110100001000011100010100000101111; end
            14'd6932 : begin out <= 64'b0010010111100000101001010000011100011101101001010010101110101100; end
            14'd6933 : begin out <= 64'b1010101110010010101010001000001110100010011110000010100001011110; end
            14'd6934 : begin out <= 64'b1010010101000010001010001010010100100011111001000010100100011100; end
            14'd6935 : begin out <= 64'b1001101111110001001010001101100110101001001000011010001101000001; end
            14'd6936 : begin out <= 64'b1010100001111000101010111110001010101011011111001010101100010110; end
            14'd6937 : begin out <= 64'b1000101010110111101001101111010100101000100001110010101100110101; end
            14'd6938 : begin out <= 64'b0010010100110011101010001110000000100100111010111010001110110010; end
            14'd6939 : begin out <= 64'b0010011100000000101001111011001000100100111110100010101011000100; end
            14'd6940 : begin out <= 64'b0010010010111100101001101111101010100000000001101010101100011000; end
            14'd6941 : begin out <= 64'b1010101111001000101001101111110010100101000010101010010110110011; end
            14'd6942 : begin out <= 64'b1010000001101100001001001100100100101010100100010010100011100010; end
            14'd6943 : begin out <= 64'b1010001011100001101010001011111000100011001001011010101101000111; end
            14'd6944 : begin out <= 64'b0010101011011111101010110011010000101011001001111010101110010111; end
            14'd6945 : begin out <= 64'b1010101010011100101010111001111010100001101100100010100001011111; end
            14'd6946 : begin out <= 64'b1010100011111000101000110100100010100010011001111010101000001111; end
            14'd6947 : begin out <= 64'b0010000011101011101001001111111010101001110101011001011010111001; end
            14'd6948 : begin out <= 64'b1010101101010111001001101011010000101010100010100010100111011101; end
            14'd6949 : begin out <= 64'b1010000111010110001001110001110110101011010111110001011010111011; end
            14'd6950 : begin out <= 64'b0010100011100111101010110111101010001011011001101010001110101110; end
            14'd6951 : begin out <= 64'b0010100101001110101010110101010100100111101001010001001101000010; end
            14'd6952 : begin out <= 64'b1010000101110000101000110011100110100011110010111010101010100101; end
            14'd6953 : begin out <= 64'b0010010001000001001010111110110100011110010111110010011111010000; end
            14'd6954 : begin out <= 64'b1010100100110100001001101011011010101010100010110010101111001101; end
            14'd6955 : begin out <= 64'b0010100110111100101001101000011000100110110101111001010010011110; end
            14'd6956 : begin out <= 64'b0010011101000111001000001001111010100010011111110010100100100000; end
            14'd6957 : begin out <= 64'b0010101100101011001010000010011110100111000100011010011000000001; end
            14'd6958 : begin out <= 64'b1010100101000001101001100110100000101010011110101010000000101101; end
            14'd6959 : begin out <= 64'b1010101110010001001010110001001000101010011111101010101011011000; end
            14'd6960 : begin out <= 64'b0010101101111011001001001111000010011110011001011010101000011101; end
            14'd6961 : begin out <= 64'b0010011111101011101000000010101000100110010101110010101010101101; end
            14'd6962 : begin out <= 64'b0010011010101010101000011100111010100110011000011010100011000011; end
            14'd6963 : begin out <= 64'b0010011111100000101001101011010100100100001110101010011110101010; end
            14'd6964 : begin out <= 64'b0010010110110001101010111011110010100110011100000010011100101110; end
            14'd6965 : begin out <= 64'b0001110010011001001001001101111110100100110100101010011010011110; end
            14'd6966 : begin out <= 64'b0010010001111000001010100111001010101001111011011010001110101010; end
            14'd6967 : begin out <= 64'b0001000101011011101010000000010000100101011010110010001010101001; end
            14'd6968 : begin out <= 64'b1010100111000010001001100111000100011111001110101001111101000101; end
            14'd6969 : begin out <= 64'b0010011010100001101001111010111010101001111011011010101010010110; end
            14'd6970 : begin out <= 64'b1010101001001100001010100000110110010001010111101010101100100001; end
            14'd6971 : begin out <= 64'b1010101101110101101010011111000110100010110000111010010100100001; end
            14'd6972 : begin out <= 64'b0010010000001110001010001100000000100101101011000010101010101101; end
            14'd6973 : begin out <= 64'b1010101000101111101010001000110110010101001100101010100110111101; end
            14'd6974 : begin out <= 64'b1010100000011100101010000100101000101000110000000010000111011110; end
            14'd6975 : begin out <= 64'b1010001101101010000111010110110000100011010000010010010011101101; end
            14'd6976 : begin out <= 64'b1010000101001000101001010111110100101001111000111010011101111111; end
            14'd6977 : begin out <= 64'b0010100000100000001011000110111000101000001101010010100111100110; end
            14'd6978 : begin out <= 64'b0010010111101101001010101100000000101000110001111010101010100110; end
            14'd6979 : begin out <= 64'b1010101111000001101000001111100100100011000000110010100000110100; end
            14'd6980 : begin out <= 64'b1001110101000110001001110110000110100110111010000010100111001011; end
            14'd6981 : begin out <= 64'b0010100000100010100110101110100100100101001100111010101111110000; end
            14'd6982 : begin out <= 64'b1010011001011110101010100011101010011100001010001010101011100010; end
            14'd6983 : begin out <= 64'b1010011111111101100110100011100110101011000100100010000110000011; end
            14'd6984 : begin out <= 64'b0001111010100101101010011111100010100010110011010010101100101110; end
            14'd6985 : begin out <= 64'b1010011101001111000011000001111110101000010001110010100000111101; end
            14'd6986 : begin out <= 64'b1010001110110011001001001110010010101001101101000001111000101011; end
            14'd6987 : begin out <= 64'b1010011111110010000110101101001000100001001111100010001111011111; end
            14'd6988 : begin out <= 64'b0010101000111111101010100110111110101010100110101001111110100000; end
            14'd6989 : begin out <= 64'b0010001100100110101010011001001110011110001011000010010111101011; end
            14'd6990 : begin out <= 64'b0010100100101111001010000110011010100101101011010010101010010000; end
            14'd6991 : begin out <= 64'b0010101110010101001010100110111100100100010001111010010111100100; end
            14'd6992 : begin out <= 64'b1010100010100010101010000101111110100000000001010010011011110110; end
            14'd6993 : begin out <= 64'b0010101101000000101001000101111010101000000100100010010110101100; end
            14'd6994 : begin out <= 64'b0010011101101100101001011010000110101000111001111010100111100001; end
            14'd6995 : begin out <= 64'b1010101101001100001010000000110110011111001011100010100001110110; end
            14'd6996 : begin out <= 64'b0010100011011101001010001110100000101001110000111010100111001001; end
            14'd6997 : begin out <= 64'b1010010110011011001010010011001100100101010101001010011000110001; end
            14'd6998 : begin out <= 64'b1010100110010111101010000010001010100101010110011010000001001011; end
            14'd6999 : begin out <= 64'b0001110000010110001010100010110100100001001001001010011011110010; end
            14'd7000 : begin out <= 64'b0010100010001010100111000101001110100011000100000010010111100101; end
            14'd7001 : begin out <= 64'b1010000111110010001001100111101100101000011010110010010111001010; end
            14'd7002 : begin out <= 64'b0010011110100110001010000010000100100010101001011010000000111111; end
            14'd7003 : begin out <= 64'b0010011101101110101001101101101110100111011110100010101111011001; end
            14'd7004 : begin out <= 64'b0010101100011001101000010001000100101011110010000010110000111000; end
            14'd7005 : begin out <= 64'b0010101001111100101010101001001010101000111010100001110000010111; end
            14'd7006 : begin out <= 64'b1010100101011000101010111111000110101011011100110010000100001101; end
            14'd7007 : begin out <= 64'b0010101000011111101010100010101010100001011100001010010001101001; end
            14'd7008 : begin out <= 64'b1010100111001000000111100011010000101011110110111010101111100101; end
            14'd7009 : begin out <= 64'b0010000101111111101000100011100000101010111110000010101110110110; end
            14'd7010 : begin out <= 64'b1010100010011101101010110111011000100011110010011010100111000111; end
            14'd7011 : begin out <= 64'b1010101010010011100100110011000010100110000011000010001111010010; end
            14'd7012 : begin out <= 64'b1010101011010111001010000000111100101001101011100010100110010111; end
            14'd7013 : begin out <= 64'b1010101101001011001000101100101100101010100001010010001111001110; end
            14'd7014 : begin out <= 64'b1010001100110101000111101010110100101011010001011010100110000011; end
            14'd7015 : begin out <= 64'b1010101110001001101010111011101110100111101010111010000010110101; end
            14'd7016 : begin out <= 64'b0010010000101001001001010010111110101011100101111001101101100101; end
            14'd7017 : begin out <= 64'b0010010100110010001010111000110010100111000010000010100001100110; end
            14'd7018 : begin out <= 64'b0010011101100101001001101111101000101010110111010010100111100100; end
            14'd7019 : begin out <= 64'b0010010000000111000111001000010110100101111111101010100011011111; end
            14'd7020 : begin out <= 64'b1001111111100011001001111100001110101000001001011010011000111001; end
            14'd7021 : begin out <= 64'b0010010000110100101010001011111100011111000010101010100011111101; end
            14'd7022 : begin out <= 64'b1010101010110110001001000101110100100111111001100010100000110110; end
            14'd7023 : begin out <= 64'b1010011001100001001000111000101000100001110100100010010001001100; end
            14'd7024 : begin out <= 64'b1010010011011001001000111011110110101000000011111010011101001101; end
            14'd7025 : begin out <= 64'b1010010101000100101010010111101110100010100001100010010101100010; end
            14'd7026 : begin out <= 64'b1010010000000011101010111010010010100110100111000001010000110011; end
            14'd7027 : begin out <= 64'b1010001001110111001001000011010110101000011001110010100001001011; end
            14'd7028 : begin out <= 64'b1010001101001111001010011000000000101001101101100010101101000110; end
            14'd7029 : begin out <= 64'b1010101100110100001010000001010000100101100000000010101010110001; end
            14'd7030 : begin out <= 64'b0001100111010010000111000011001010101001111111111010101100110100; end
            14'd7031 : begin out <= 64'b0001000010001110001001100100100110010011001111110010001001110000; end
            14'd7032 : begin out <= 64'b1010100000101001001010101100111000101001101110000001111011000010; end
            14'd7033 : begin out <= 64'b1010001110000101101001111110101000011000010010110001010000001000; end
            14'd7034 : begin out <= 64'b0010011000111001101011000001110100100001110111010010101101110101; end
            14'd7035 : begin out <= 64'b0010101011010110001010101010010110010010000011111010100110101010; end
            14'd7036 : begin out <= 64'b0010100001000011001010010110111100100011101011111010100000101001; end
            14'd7037 : begin out <= 64'b1010100110111101101010111010011000100100001100010010101110111111; end
            14'd7038 : begin out <= 64'b0010001101011010000110111001100010100010010100101010010001111010; end
            14'd7039 : begin out <= 64'b0010010101001101101010000111010110101001111000110010100000101110; end
            14'd7040 : begin out <= 64'b1010100101110110100111100000110100101011011110011010100001111010; end
            14'd7041 : begin out <= 64'b1001011101011101001010010111101010100000111111011001111110001110; end
            14'd7042 : begin out <= 64'b0010011000000110101001000111011010101001111111001010000101001101; end
            14'd7043 : begin out <= 64'b1010100101100100001010111101001000101000111101010010110000110101; end
            14'd7044 : begin out <= 64'b1000011111111000101010111100111010101000010111000010101000101000; end
            14'd7045 : begin out <= 64'b0010011111100101101010001001000010101011011110101010101101010110; end
            14'd7046 : begin out <= 64'b1001111000111000001001101111101100101000100000011010101001010111; end
            14'd7047 : begin out <= 64'b1001110101010011001001001000011000101000011010110010001111010001; end
            14'd7048 : begin out <= 64'b1010100111101110001010001011110010100001110001110010100010000111; end
            14'd7049 : begin out <= 64'b0010110000001001101010011010010010010010101010000001110110001000; end
            14'd7050 : begin out <= 64'b1010010101000111001010010010111100101010111010110001110111100110; end
            14'd7051 : begin out <= 64'b1010100100111000000011100000111000100110011111101010010101010000; end
            14'd7052 : begin out <= 64'b1010101110101000000111110101010010101010010010110010100001111011; end
            14'd7053 : begin out <= 64'b1010000110110011001000011000111000100110001000101010001101101011; end
            14'd7054 : begin out <= 64'b0010001100110101101001111111001100100110011101110010010000101100; end
            14'd7055 : begin out <= 64'b0001111100100111101010011111001100101001110011100010001001001111; end
            14'd7056 : begin out <= 64'b0010100000100101101010100101111010101010000101010010100001000010; end
            14'd7057 : begin out <= 64'b0001100111000101101010010001111010011000001010011010100101010011; end
            14'd7058 : begin out <= 64'b1010100000011101001010010000011010100011111011101010101010010010; end
            14'd7059 : begin out <= 64'b0010000100001010101010011111111110101010000000110010101010011110; end
            14'd7060 : begin out <= 64'b0010010010000110101001111110001010011101011000100010011110000110; end
            14'd7061 : begin out <= 64'b0010101111001010101001111001111110100000100010110001100100010110; end
            14'd7062 : begin out <= 64'b1010101001011110001001000010001110011010001111100001011101101100; end
            14'd7063 : begin out <= 64'b0010100011101010101010011110001010100100001001110001101000010010; end
            14'd7064 : begin out <= 64'b1010011111111001101010000101110110101000101011011010100101100110; end
            14'd7065 : begin out <= 64'b0010001101111100001010011010100110011110010011101010100111100000; end
            14'd7066 : begin out <= 64'b1010011010100011001001010000110010101011010010001010010001110110; end
            14'd7067 : begin out <= 64'b0010011101001101001010110111010010101010010010010001110010000110; end
            14'd7068 : begin out <= 64'b0001010000100101101010010010111010101011101001100010101001001100; end
            14'd7069 : begin out <= 64'b0001111101111001000010101101011000100111110100100001000111000100; end
            14'd7070 : begin out <= 64'b0010010000000110001010111100000100000101011110001010010010000000; end
            14'd7071 : begin out <= 64'b1010101010110101001010001011100110100011000100011010101110000110; end
            14'd7072 : begin out <= 64'b1010011101110111101010010010001110101010100000010010001100010011; end
            14'd7073 : begin out <= 64'b0001110010011000001000010001010010100100110110101010010010010100; end
            14'd7074 : begin out <= 64'b1010101000101011101000010101100010101000100101010010101100010100; end
            14'd7075 : begin out <= 64'b0010001000110110101010001001010000011010110100001010000111111100; end
            14'd7076 : begin out <= 64'b0010101110011111001010101100111110100100110011011010011110110100; end
            14'd7077 : begin out <= 64'b1010010111001111001010011100110010100000100000110010100000100000; end
            14'd7078 : begin out <= 64'b0010100000101010001010000000101000100111001111100010011101000110; end
            14'd7079 : begin out <= 64'b0010001111101111101011000100101100101000001100101010100000100101; end
            14'd7080 : begin out <= 64'b0010101110111000101010011100010100100111000001000010100101110111; end
            14'd7081 : begin out <= 64'b0010100101100100100110011110000010101000001111110010000011011111; end
            14'd7082 : begin out <= 64'b1010010101110001101001111011000100101010001110100010100100111111; end
            14'd7083 : begin out <= 64'b0010010100110011101011000011010010100101110000000010100001001111; end
            14'd7084 : begin out <= 64'b0001111001000011001000001110111110101000101111010001101111111100; end
            14'd7085 : begin out <= 64'b0010011000111100001010101001100110100110101101010010010001110000; end
            14'd7086 : begin out <= 64'b1001111110100000000111001101100100101001011111011010011100111100; end
            14'd7087 : begin out <= 64'b0010100111011000000101110100111010100111111101001010101001001001; end
            14'd7088 : begin out <= 64'b1010101011011001000110110111000000101000110010001010011100011100; end
            14'd7089 : begin out <= 64'b1010100011000100101001110101010110101001010100110010100101111101; end
            14'd7090 : begin out <= 64'b0010100011110101101010001000111110101011011110111010000001101000; end
            14'd7091 : begin out <= 64'b0010101010011101101010011000100010100100101110010010001001101101; end
            14'd7092 : begin out <= 64'b0010101010111011101010110011011010101011000111111010100010001011; end
            14'd7093 : begin out <= 64'b0010001000001010101000110110101110100101100010010010101101000101; end
            14'd7094 : begin out <= 64'b1010100001111001001010011111101000100010010101100010000010011111; end
            14'd7095 : begin out <= 64'b0010100000001110101001100111100110100100011011111010100100111100; end
            14'd7096 : begin out <= 64'b1010010111100111101000100111110000101011011001111010001010111111; end
            14'd7097 : begin out <= 64'b0010001111101110101000011100111010100001011100111010100010001101; end
            14'd7098 : begin out <= 64'b1010100100000101101010000011100110101010111000001010100111000010; end
            14'd7099 : begin out <= 64'b1010011011010011001001111011000010100111000000010010100000010011; end
            14'd7100 : begin out <= 64'b1010011011101101101010011100110110101011100000111010010100101010; end
            14'd7101 : begin out <= 64'b0001011000011101100111100001101000101000111010011001110010011101; end
            14'd7102 : begin out <= 64'b0010010010100110001001011100000010101010001101111010011100010010; end
            14'd7103 : begin out <= 64'b0001110011000001000110010100100000100100011001000001111100001101; end
            14'd7104 : begin out <= 64'b0010101101010101001000111001011000100100101101111010101010010111; end
            14'd7105 : begin out <= 64'b0010101010111100101010011100100110100101101000011010110000000010; end
            14'd7106 : begin out <= 64'b1010100011100101101010011000010000100001111011111010001101010001; end
            14'd7107 : begin out <= 64'b0010101010000111001001011010100100100110010101001010010110001100; end
            14'd7108 : begin out <= 64'b0010011111100100101001101011101010100101010001111010011101011110; end
            14'd7109 : begin out <= 64'b1010100001111010001001101001010100101010001100101001100000110001; end
            14'd7110 : begin out <= 64'b0010100101111101001001001111010000100100100010110010010011010100; end
            14'd7111 : begin out <= 64'b0000100111010010001010110011001010101000111110011010101101011100; end
            14'd7112 : begin out <= 64'b1001111101010011101010100001001000101010010011100010000100100111; end
            14'd7113 : begin out <= 64'b1010101101110100101001111111010010100110000000101010100101001111; end
            14'd7114 : begin out <= 64'b1010110000000100000110011010010100101010101110010010011100110000; end
            14'd7115 : begin out <= 64'b1010101100001111001000000011010110100001101111001001100101111010; end
            14'd7116 : begin out <= 64'b0010100000011110001001111010000010101010010101010001101000100011; end
            14'd7117 : begin out <= 64'b1010000000101111101010110000010110100101001010010010011110000110; end
            14'd7118 : begin out <= 64'b1010101100010011001000110001000100101001011000001010100011011010; end
            14'd7119 : begin out <= 64'b0010010001110110001001001010010000100111100111000010100011001101; end
            14'd7120 : begin out <= 64'b1010100100100011001010010110100100100111001000011001111101100100; end
            14'd7121 : begin out <= 64'b0010001101000001001010101111001000101010011001010010100101010101; end
            14'd7122 : begin out <= 64'b0010000111001101001001000001110110101001110001010010010100100100; end
            14'd7123 : begin out <= 64'b0010010100111100101000101110110010101001100111101010101111111110; end
            14'd7124 : begin out <= 64'b1010011010100001101010001000011000011001010000100010001011001101; end
            14'd7125 : begin out <= 64'b0010011001110110001000100001110100101000010100010010101000000100; end
            14'd7126 : begin out <= 64'b1010000100110010101010010010100100100001101111011010100000000010; end
            14'd7127 : begin out <= 64'b0010101000111000101010000100000010101000001111101010101110101111; end
            14'd7128 : begin out <= 64'b0010100111010011001010000111100100101010101001011010010111011001; end
            14'd7129 : begin out <= 64'b1001011100101101001000011010100100101001101111100010010010011000; end
            14'd7130 : begin out <= 64'b0010101011010010001001000111011110101001011100001010100001010111; end
            14'd7131 : begin out <= 64'b1010101000000001001000100011000100100000110000000010101101011100; end
            14'd7132 : begin out <= 64'b1010101000001100001001011010111000101000011000101010100000010000; end
            14'd7133 : begin out <= 64'b0010010110111111000011001101101000101010100011011001010011110100; end
            14'd7134 : begin out <= 64'b0010100110111000101001000100010100101011011100101001010101000000; end
            14'd7135 : begin out <= 64'b0010101001101010001010010101000110100110001100001010011001010100; end
            14'd7136 : begin out <= 64'b0010010000000111101010000000000100100101010101011010100001011101; end
            14'd7137 : begin out <= 64'b0010011100101010001010101000000100101011001011100010100111001110; end
            14'd7138 : begin out <= 64'b0001111101011110001010111010011000101000100000010010000100010100; end
            14'd7139 : begin out <= 64'b1010101100101110001000000101011100011110011101100010101011001110; end
            14'd7140 : begin out <= 64'b1010101101110111001010110110110000101000001111000010000000000001; end
            14'd7141 : begin out <= 64'b1010100000000110001010111001001100101011111101011010010110101110; end
            14'd7142 : begin out <= 64'b1001111010101001001000010111110100100010011000011010011111100001; end
            14'd7143 : begin out <= 64'b0010001110100111000111110101001000100001011000101010100110110101; end
            14'd7144 : begin out <= 64'b1010010001011100100111001010001100101010110011001010000010110100; end
            14'd7145 : begin out <= 64'b1010101010010001001010100001010110100011010100001010001111100011; end
            14'd7146 : begin out <= 64'b1010010010000000101010110110011010100101001110001010101100011101; end
            14'd7147 : begin out <= 64'b0010001100000001101010110011101010101010010111011010101110000000; end
            14'd7148 : begin out <= 64'b0001011001111001001001111100001110101000100101111010101101001111; end
            14'd7149 : begin out <= 64'b0010101101010110101001000101011100101001110001111010011110011100; end
            14'd7150 : begin out <= 64'b0001001100100011000101011101001010101000101010100010100000111100; end
            14'd7151 : begin out <= 64'b1010101000000111001011000101000110100110011001110010011101001011; end
            14'd7152 : begin out <= 64'b0010100100111010100111011010011000101011101001001010010010011011; end
            14'd7153 : begin out <= 64'b1001100011101000001010011110011110100110000000010010001111010101; end
            14'd7154 : begin out <= 64'b1010011010100101001010110010001010101011010111110010100010110000; end
            14'd7155 : begin out <= 64'b1010001001011011101010101111010010101000001100101010101110011001; end
            14'd7156 : begin out <= 64'b1010010110011100001001010011100110010011010110010010100001110100; end
            14'd7157 : begin out <= 64'b1010010100111110001001100011001010101000000001100001111111010101; end
            14'd7158 : begin out <= 64'b0010100100011110101010101011101000011011001011111001111111111100; end
            14'd7159 : begin out <= 64'b1010010110011110001010001011011000101001111011010010100101000111; end
            14'd7160 : begin out <= 64'b1010100011010100101000111110100100100101100010111001101111101000; end
            14'd7161 : begin out <= 64'b0010100111101001001010101110110000101011111111111010011111101101; end
            14'd7162 : begin out <= 64'b1010100001001111101010110001000100100110000000111010100110101010; end
            14'd7163 : begin out <= 64'b0010100001100111100111101111001110100101101111111010101101000011; end
            14'd7164 : begin out <= 64'b0010100001011100001010010011101000100110011100000010101101111001; end
            14'd7165 : begin out <= 64'b1010010100100110101010111001001010011111000011011010101010100110; end
            14'd7166 : begin out <= 64'b1010100110111001001010011101001110101010111001110010011101000111; end
            14'd7167 : begin out <= 64'b0010101110101111001000110111100100100000110110101001111110101011; end
            14'd7168 : begin out <= 64'b1010101010101011001001110101111100101011110110000010010100101001; end
            14'd7169 : begin out <= 64'b0010010111111110001000000100110110100001100111000010101010000001; end
            14'd7170 : begin out <= 64'b1001110011000001100110011000011000100000011111101001100011111110; end
            14'd7171 : begin out <= 64'b0010001010100100101000100010100000101001110000101010010110110100; end
            14'd7172 : begin out <= 64'b0010010111011011001010011110100010100010110010101010100001100001; end
            14'd7173 : begin out <= 64'b1010101001001101100111011111010010100000101110001010010111011101; end
            14'd7174 : begin out <= 64'b0010100001000111001010010001010000100110110010011010101110111100; end
            14'd7175 : begin out <= 64'b1010101001100000001010101000011100100100010110100010011101011101; end
            14'd7176 : begin out <= 64'b1010001011111110101010101110001000011110000101011010101000011100; end
            14'd7177 : begin out <= 64'b0010100000010010101010100101100100101011011010000001100110110100; end
            14'd7178 : begin out <= 64'b0010101001110001001010110110010010101001011000011010001100011001; end
            14'd7179 : begin out <= 64'b1010100101010101001010011000000010100100110110101010010100110001; end
            14'd7180 : begin out <= 64'b0010001110111101101000111011010000100101010001101010101111101100; end
            14'd7181 : begin out <= 64'b1010000010000111101010001111110110100110010010010010101000011000; end
            14'd7182 : begin out <= 64'b1010100100001001001010100000001110100010011101101010100111110000; end
            14'd7183 : begin out <= 64'b1001101111101001101010100101110000100011110001011010011011000100; end
            14'd7184 : begin out <= 64'b1010010010000100000101110110010110100101010001001010010010100011; end
            14'd7185 : begin out <= 64'b0010100110010010001010011100001000100100101100111010010101110010; end
            14'd7186 : begin out <= 64'b0010100110001010101010000100101110100111001011100010011110001001; end
            14'd7187 : begin out <= 64'b0010000010000010001001111000111110100111110001110010100011000101; end
            14'd7188 : begin out <= 64'b1010100111111011100111010111110110100110111000110010011111111111; end
            14'd7189 : begin out <= 64'b1001010110110000101000101110100100101000000000011010001100011100; end
            14'd7190 : begin out <= 64'b1010001001010111001000001101100110100000011000010010001000000001; end
            14'd7191 : begin out <= 64'b0010101000101110101010111011101000101010111011001001111111101010; end
            14'd7192 : begin out <= 64'b1010101101100111001010010110100000101010001111011010100110001111; end
            14'd7193 : begin out <= 64'b1010010101110000101010010101111110101010000001010010101101101011; end
            14'd7194 : begin out <= 64'b1010101101111011101010110111101100100101001111101010100011111000; end
            14'd7195 : begin out <= 64'b1010101001011100101000010101110110010101011000001001111111011101; end
            14'd7196 : begin out <= 64'b1010100110100111101010001010011100100101110110110010010101010011; end
            14'd7197 : begin out <= 64'b1010101100100011101010111001101100101011111001011001011101111100; end
            14'd7198 : begin out <= 64'b1010100010101101001001000001110110011100110111011010000010111111; end
            14'd7199 : begin out <= 64'b0010011101101011101010100010100010011000001100111010110000010101; end
            14'd7200 : begin out <= 64'b1010101011011000101010011110000100100100010100000010100111000110; end
            14'd7201 : begin out <= 64'b0001111010110110101010111100000110100010000011100010100111110000; end
            14'd7202 : begin out <= 64'b1010100101111111001001010011101100101011011100001010101010010100; end
            14'd7203 : begin out <= 64'b0010101000100011101010011111101110100110000111011010011010011000; end
            14'd7204 : begin out <= 64'b0010010111001110001010011001101110100110111111111010100010110000; end
            14'd7205 : begin out <= 64'b0010101110110011101010100000011100101010111011011010100110010101; end
            14'd7206 : begin out <= 64'b1010000111100001101010011100000100101010011001101010100011111111; end
            14'd7207 : begin out <= 64'b1010010001100000001010111100101110101010011001100010011100110011; end
            14'd7208 : begin out <= 64'b0010000001001111101010001000010100101001010101110001101100111110; end
            14'd7209 : begin out <= 64'b1010000110010011101001101111011000100111110010000010010010001110; end
            14'd7210 : begin out <= 64'b0010010101010110001010110000110010101010011111110010101000101110; end
            14'd7211 : begin out <= 64'b0010100110100001001010010010101110100100011010010010101110101001; end
            14'd7212 : begin out <= 64'b1001111110000000101001000111111010100111101010110010101111011101; end
            14'd7213 : begin out <= 64'b0010010000001010101001000100111000101001011011101001111111110010; end
            14'd7214 : begin out <= 64'b0010110000010011101000100011111000101000100011000010010111101110; end
            14'd7215 : begin out <= 64'b0010101010100011001010010011111100101000101010010010100000111011; end
            14'd7216 : begin out <= 64'b0010101110011000100110110011100000101010001001000010010010011010; end
            14'd7217 : begin out <= 64'b0010001011111100101010111000110000101010111101100010100100011001; end
            14'd7218 : begin out <= 64'b0001011100011100000111111101100110011101001010110010100100000010; end
            14'd7219 : begin out <= 64'b1010000000010110001000111100101110101010000100011010101001101101; end
            14'd7220 : begin out <= 64'b0010101000000100000111010101010100101011010001111010101100011111; end
            14'd7221 : begin out <= 64'b1001111000100101001010100011000000100100001100010010101100100101; end
            14'd7222 : begin out <= 64'b1010001011001001101001110111001000100110000011010010101001001000; end
            14'd7223 : begin out <= 64'b0010100111100010101001010000001100101011101010011010011111000110; end
            14'd7224 : begin out <= 64'b1010100011011001001010001011100110101011111011010010100001101010; end
            14'd7225 : begin out <= 64'b0010001111011100001001000011000110011010110100001010001000101001; end
            14'd7226 : begin out <= 64'b0010001111000010000111011001010000101000001100011010101000000010; end
            14'd7227 : begin out <= 64'b0010001000000010001010111001101110100000110000100010010010110000; end
            14'd7228 : begin out <= 64'b1010011010100111001010001000110110101001001001011010110000100110; end
            14'd7229 : begin out <= 64'b0010000110100001001001100111101000101001001000010010010101001000; end
            14'd7230 : begin out <= 64'b0010011110011100001010111001010100101010010001001010010100101001; end
            14'd7231 : begin out <= 64'b0010011010000110001010100110110100100100110110010010011011001010; end
            14'd7232 : begin out <= 64'b1010010101111100001001111010101000101000101101011010100101001101; end
            14'd7233 : begin out <= 64'b1010101001110110001010100101100000101011000111011001110011100111; end
            14'd7234 : begin out <= 64'b0010010101001000101010100100111010100011010110000010011100101111; end
            14'd7235 : begin out <= 64'b0010001011100010101010000111000100011000000111100010100011110011; end
            14'd7236 : begin out <= 64'b1010100101101000101001101100101000011100100011100010010000010110; end
            14'd7237 : begin out <= 64'b0001001001111010001010001011000000101001101010011010000011110001; end
            14'd7238 : begin out <= 64'b0010100110001110000100110000100010100100110110100010100000000111; end
            14'd7239 : begin out <= 64'b0000110001101111100110001101100000011010010100010010101001101100; end
            14'd7240 : begin out <= 64'b1010101000010110100111001110100100011000111010010001101100100111; end
            14'd7241 : begin out <= 64'b1010010011100100000110000111001010101011001010001010101010111101; end
            14'd7242 : begin out <= 64'b1001110110000101101010010101111010100010111100010010101100001000; end
            14'd7243 : begin out <= 64'b0010100100110010101010010001000110101011000110011001011101001000; end
            14'd7244 : begin out <= 64'b0001010100101011000111111101110000100101010101100010100111110010; end
            14'd7245 : begin out <= 64'b1010100101110001100110010000111000100110100100100010011100000111; end
            14'd7246 : begin out <= 64'b1010100001001001001001111101011110101000100100010010100100001110; end
            14'd7247 : begin out <= 64'b1010010001011110101010111011000110100101100101111010100000110111; end
            14'd7248 : begin out <= 64'b0001101100001101101001001100010100101010100100010010000100101001; end
            14'd7249 : begin out <= 64'b0010010000111100001001000111000100101010101010101010101110110101; end
            14'd7250 : begin out <= 64'b0010011011010001101000101000000110100010100101011010101110010011; end
            14'd7251 : begin out <= 64'b1010001101011010101001101110110000101001111101010010011101001100; end
            14'd7252 : begin out <= 64'b1010011011011000001010001000111110101000011101111010011001111100; end
            14'd7253 : begin out <= 64'b0010100101100101101010110010100100101010001101110010100101000000; end
            14'd7254 : begin out <= 64'b1010001001101100001010001101100010011111000001000010101011001001; end
            14'd7255 : begin out <= 64'b1010101100100010101001111100111000100111110111111010100110000000; end
            14'd7256 : begin out <= 64'b0010000001000001101010001010101000100110111000101010000000110011; end
            14'd7257 : begin out <= 64'b1010010100111101101010000111010010100001110010010010100001110001; end
            14'd7258 : begin out <= 64'b0010100010010001001000100100001000011110010111100010101111001110; end
            14'd7259 : begin out <= 64'b1010100111000010101010100110010010101001000000010010011101100100; end
            14'd7260 : begin out <= 64'b0010010100111000001010110000001100101000010111011001100101101011; end
            14'd7261 : begin out <= 64'b1010011010101101101010100111010010100011100101011010101101010101; end
            14'd7262 : begin out <= 64'b1010100011011110101010100110110000101010011000101010101011101101; end
            14'd7263 : begin out <= 64'b1010100010001101001000011111111100011110100110000010011100011000; end
            14'd7264 : begin out <= 64'b1010011101110110101010110010101100011000101000111010001001001001; end
            14'd7265 : begin out <= 64'b0001111111000010001001110011111110100101110001010010100011111111; end
            14'd7266 : begin out <= 64'b0010101110110111001000111001010100100100111101001010011011011000; end
            14'd7267 : begin out <= 64'b1001111111111110001000000000011110011101110100101010011001001010; end
            14'd7268 : begin out <= 64'b0010101100000010001001011000100000100001001111111010100110000100; end
            14'd7269 : begin out <= 64'b1010100010001001001001010101111000101011101011000010100101110000; end
            14'd7270 : begin out <= 64'b1010100101000010001010011111101010101000101110101010011010101100; end
            14'd7271 : begin out <= 64'b0010000011001001101001111000101110100010010111100010010111011100; end
            14'd7272 : begin out <= 64'b1010100101010101101010000101010000100010101001101010101001101111; end
            14'd7273 : begin out <= 64'b0010001101101100101010001011100100101010110101101010100001101010; end
            14'd7274 : begin out <= 64'b0010000010000011101001010101101110101000011011011001101001001000; end
            14'd7275 : begin out <= 64'b0010101000001011001010011111000010101010101001110010100101000000; end
            14'd7276 : begin out <= 64'b1010100010000011001001101100000000101011101011101010010111101100; end
            14'd7277 : begin out <= 64'b1010101000110100101010111111011000100101000111001010000100010110; end
            14'd7278 : begin out <= 64'b0010101001010100001010001010111110101001111011010010100101011011; end
            14'd7279 : begin out <= 64'b1010101110001110001001000100001100101001000001100010110000001011; end
            14'd7280 : begin out <= 64'b1010001010111010101000100010001000011101011101010001110101101110; end
            14'd7281 : begin out <= 64'b0010101110010011101001111010010000101011010011100010100000000111; end
            14'd7282 : begin out <= 64'b1010101101110010000110001001111010011000011011010010101010101001; end
            14'd7283 : begin out <= 64'b1010101011011011101010000100111110101011001001001010011010000101; end
            14'd7284 : begin out <= 64'b1010010111100011001010100010100100100010111100010001111101111111; end
            14'd7285 : begin out <= 64'b1001101000001001101010111000001000101001111010100010000100011100; end
            14'd7286 : begin out <= 64'b1001011000110000001001000101000100100110000010001010101001110100; end
            14'd7287 : begin out <= 64'b0010100110111110101010000000101010101000011010100010100011101111; end
            14'd7288 : begin out <= 64'b0010001111001010001010011100101010101010010011011010100100100000; end
            14'd7289 : begin out <= 64'b1010101110011001001010101000011110100100100000111010100000010100; end
            14'd7290 : begin out <= 64'b0010100000101110101010010000110100100101100101111010100011001001; end
            14'd7291 : begin out <= 64'b0010101010011011001010100001110000100000101101000001000010000110; end
            14'd7292 : begin out <= 64'b0010011101010010101010111110110010100110001101101010100000111110; end
            14'd7293 : begin out <= 64'b0010100001001000101000110110001000101000010110000010100111100000; end
            14'd7294 : begin out <= 64'b0010101011011110000101000010111110101011000101001010001101001001; end
            14'd7295 : begin out <= 64'b0010011010010101000110101111110000100010001000101010100100010000; end
            14'd7296 : begin out <= 64'b1010100010101100000101010010110100101011100000011010010100011011; end
            14'd7297 : begin out <= 64'b1010101001010001100111010001010000100100001011101010000001011000; end
            14'd7298 : begin out <= 64'b1001001110110011100110001111100000101000111011001010100111111001; end
            14'd7299 : begin out <= 64'b0001101101101010101000010011101100101001010100011010010101100010; end
            14'd7300 : begin out <= 64'b0010010000010011100111000011000100101000010100000010001000010011; end
            14'd7301 : begin out <= 64'b0010101001001111001001111110010100100100101011001010101101010001; end
            14'd7302 : begin out <= 64'b0010100100110110001001110100011110100111111111000010011110000110; end
            14'd7303 : begin out <= 64'b0001111001000000101001011100111100101010001101101010001010101001; end
            14'd7304 : begin out <= 64'b0010100010101000101000100110011110101010111111010010100110111010; end
            14'd7305 : begin out <= 64'b0010000111100000001010111011100010100111010100110010101011111001; end
            14'd7306 : begin out <= 64'b0010011101000000101001110100011100100001010000110010100100100011; end
            14'd7307 : begin out <= 64'b1010000010110111101010010000000110100111011001000010101110100000; end
            14'd7308 : begin out <= 64'b0010000100101101001010100111111010101010100011110010101000100001; end
            14'd7309 : begin out <= 64'b1010101100010111100110001100000010100110001000110010101000111111; end
            14'd7310 : begin out <= 64'b0010100000111111001010100010011110100101000010110010100001001001; end
            14'd7311 : begin out <= 64'b1010100110111111100100100100111110100100100110111010010111001001; end
            14'd7312 : begin out <= 64'b0001111111011001101010110100110110101001011111001001010100100011; end
            14'd7313 : begin out <= 64'b1010011100000111001010110001010100100001010011010010101111011011; end
            14'd7314 : begin out <= 64'b0010010100101001101010011100010000101000110010101010101000110010; end
            14'd7315 : begin out <= 64'b0010010101001001101000111100110000100010101011000001110001101000; end
            14'd7316 : begin out <= 64'b1010011110100011101010100110110000100010001001010010101100010010; end
            14'd7317 : begin out <= 64'b0010100010110100101000011000110100101000101011001010001110111111; end
            14'd7318 : begin out <= 64'b0001001000111100001001110111111010101010110100110010101011010010; end
            14'd7319 : begin out <= 64'b0010100001010110101010100100010010101001001101011010010000000110; end
            14'd7320 : begin out <= 64'b1010100101000101001001001110100010101000111110110010101100100111; end
            14'd7321 : begin out <= 64'b1010011001110001000111000110110010100100101111110001111011110001; end
            14'd7322 : begin out <= 64'b0010001100000011101001100011110100101001010001011010011010111000; end
            14'd7323 : begin out <= 64'b0010011101110011000100011101010100011111111110010010000111010100; end
            14'd7324 : begin out <= 64'b0010010101010001100111010001101110101001101101010010101001010000; end
            14'd7325 : begin out <= 64'b0001110100111011001010010111011010101010101100100010011011010011; end
            14'd7326 : begin out <= 64'b1010101000101000100110100100000000100101100100110010101101010110; end
            14'd7327 : begin out <= 64'b0010010011000101001010001010011110101010101010101010100001000011; end
            14'd7328 : begin out <= 64'b0001111010010011001001010001100000011001111110010010100010101011; end
            14'd7329 : begin out <= 64'b1001100111001111001010111010010010101001001110001010011100101101; end
            14'd7330 : begin out <= 64'b0010100011101100101010010110000100100110011001011001001010110000; end
            14'd7331 : begin out <= 64'b1010110000010110001010000011001110100101101111110010001101100111; end
            14'd7332 : begin out <= 64'b0010100001010110100110001000000100100110000010110010001111011100; end
            14'd7333 : begin out <= 64'b1010010100000100001010010111100000101000110000001010100010000110; end
            14'd7334 : begin out <= 64'b1010100001010001001001011111000000100110100010001010101000000101; end
            14'd7335 : begin out <= 64'b0010010000111101100111111000010010101000111000001010010101101111; end
            14'd7336 : begin out <= 64'b0001111101001011101010011101011100100111011011001010101000010110; end
            14'd7337 : begin out <= 64'b0010101010001011001000100100001100101000000001000010100001111010; end
            14'd7338 : begin out <= 64'b1001110001000110101000111011101010001011100100100010010111111000; end
            14'd7339 : begin out <= 64'b0010100010100101101001010001111100101001001000001000110000000011; end
            14'd7340 : begin out <= 64'b1010011000101100001010111001011100101010100011010010101001110101; end
            14'd7341 : begin out <= 64'b0010100001001011101010100110111010100111111100101010011101110110; end
            14'd7342 : begin out <= 64'b0010011010111100101001101001110000101010111001110010101010000011; end
            14'd7343 : begin out <= 64'b0010100011100011101001111100001110101010001000010010101001101000; end
            14'd7344 : begin out <= 64'b1010000000000110100010001011111110101000011110011001001000010110; end
            14'd7345 : begin out <= 64'b1010100110111011001010011010010110100110000001001010001000001001; end
            14'd7346 : begin out <= 64'b1010100100100100101001010010010000101001110001110010100100100100; end
            14'd7347 : begin out <= 64'b1010110000010010001010011101000000100110011101111010010000101000; end
            14'd7348 : begin out <= 64'b0001100111011110101010010101100110100000100100000010011111101110; end
            14'd7349 : begin out <= 64'b0001111001101011101010111000101110101001001010101010011101011011; end
            14'd7350 : begin out <= 64'b1010100100100111101010010110011000101011100101100010011101011110; end
            14'd7351 : begin out <= 64'b0010011100011101101010011001011100101010100100110001110001101110; end
            14'd7352 : begin out <= 64'b1010011100101001101001111011000010101000010010100001111110001111; end
            14'd7353 : begin out <= 64'b1010010011111111101001101011000010101011111010010010100001000110; end
            14'd7354 : begin out <= 64'b1010101001010100001010011011001010100011101000001010000011100101; end
            14'd7355 : begin out <= 64'b0010101111110011101010000011110010100110111100001010011011011011; end
            14'd7356 : begin out <= 64'b1010100110001110001010111111101100100011001011011010101100000011; end
            14'd7357 : begin out <= 64'b1010101101000100001010111110110010101001101100010001011000100010; end
            14'd7358 : begin out <= 64'b0010011010011001101001011001000110100001010001001010011011000100; end
            14'd7359 : begin out <= 64'b0010010100011110101010010010111100100111010011001010100010111011; end
            14'd7360 : begin out <= 64'b1001110101110110101001001101001110101011000011011010010111101000; end
            14'd7361 : begin out <= 64'b0010100100000101101010111110011100101010001100101010100001001001; end
            14'd7362 : begin out <= 64'b0010010101111000001000111001101000101001010000101001110000101001; end
            14'd7363 : begin out <= 64'b1010100011010001101010101101011000101010010111110010000111111001; end
            14'd7364 : begin out <= 64'b0010100100100000001000010011000010100111000011111010101110111000; end
            14'd7365 : begin out <= 64'b1010100101100101001010001000101010101000110011100010000011010100; end
            14'd7366 : begin out <= 64'b0001100110011100001010111011000010100110001011000010011010100010; end
            14'd7367 : begin out <= 64'b0010101001110010001010110100111010100000100111101010101101010001; end
            14'd7368 : begin out <= 64'b0010101001001011001010011100101000101011100110001010011011100010; end
            14'd7369 : begin out <= 64'b0010011111110010000111110111110010000010110100011010100110110100; end
            14'd7370 : begin out <= 64'b1010100001101001101010000000001110101010010110000001110010011001; end
            14'd7371 : begin out <= 64'b1010010101111000001001111000100000100101111010001010101110100100; end
            14'd7372 : begin out <= 64'b1010000010010100101010001110010110100101111111001010100101101101; end
            14'd7373 : begin out <= 64'b0010000001101011001010011010011010101011100010110010101111010110; end
            14'd7374 : begin out <= 64'b0010101010111010001001110001110000101001101011111010010101111010; end
            14'd7375 : begin out <= 64'b0010101110011110101010111001010000100111000000000010001010111101; end
            14'd7376 : begin out <= 64'b0010010000101100101010001110101010100011100010110010011111111101; end
            14'd7377 : begin out <= 64'b0010000010001101101010000101000010100010111001111010000001110011; end
            14'd7378 : begin out <= 64'b1010100000000111101001010100001000101000001111000010100011010001; end
            14'd7379 : begin out <= 64'b1010000010010110100101110010011110011000100011000010011101101110; end
            14'd7380 : begin out <= 64'b0010010010101111101010011111011010100100100101101001111110100111; end
            14'd7381 : begin out <= 64'b0010100001011001001010001110000100100110111010001010011000110110; end
            14'd7382 : begin out <= 64'b1010101000011110001010101101111100001111010011101010011011110101; end
            14'd7383 : begin out <= 64'b0010011100100110001000100101000110101011110001110010001000010010; end
            14'd7384 : begin out <= 64'b0010100000001000001010010000111100011000101100101010101100010101; end
            14'd7385 : begin out <= 64'b0001100100001110001010110010000010101010101100110010100011100110; end
            14'd7386 : begin out <= 64'b0010010011110100000111111010111110100010011111011010100001010101; end
            14'd7387 : begin out <= 64'b0010100110000010101000110100100000101010100011100010101110111010; end
            14'd7388 : begin out <= 64'b1010101100101111001010111100101110100100011011011010101010111100; end
            14'd7389 : begin out <= 64'b1010101100010001001010111100010010011111011011110010101010000111; end
            14'd7390 : begin out <= 64'b1010100100011100101000000011011110101010011000010010100011011011; end
            14'd7391 : begin out <= 64'b0010100001010000101001110010000100100101011100000010010001100001; end
            14'd7392 : begin out <= 64'b1010010111110011101010001101010110100100101101000010011001001010; end
            14'd7393 : begin out <= 64'b1010100100010011000100001100101010101000110101001001011101011110; end
            14'd7394 : begin out <= 64'b1010010001110111001010101000000010100101101111110010001101110110; end
            14'd7395 : begin out <= 64'b0010100101001011101001100011011010101011101101010010011101111101; end
            14'd7396 : begin out <= 64'b1010100101100011101010111010110000100101110000000010101011010111; end
            14'd7397 : begin out <= 64'b1010100100110000001010010000001100101010001001101010011011011111; end
            14'd7398 : begin out <= 64'b1010010000100011101001100000000110101010101111100010101100111001; end
            14'd7399 : begin out <= 64'b1010100111101111001010101010000110100000110011101010100010110001; end
            14'd7400 : begin out <= 64'b1010000000110001101000001101000010101011011010010001101000100111; end
            14'd7401 : begin out <= 64'b0010100000110111001010110000100110101010000111001001100010110111; end
            14'd7402 : begin out <= 64'b0010101011110110101000011011011100101010111001000010100000001001; end
            14'd7403 : begin out <= 64'b1010100001000110001010010010101010100001111101110010101111010101; end
            14'd7404 : begin out <= 64'b1010101001101110001001000010111110011100010001000010100010111100; end
            14'd7405 : begin out <= 64'b0010001110101110101010101000100010101001101111001010100100000111; end
            14'd7406 : begin out <= 64'b1010001010011110001010000100101110010110011111100010000111011110; end
            14'd7407 : begin out <= 64'b0010101000101111101000011000011000101010110101101010000100110001; end
            14'd7408 : begin out <= 64'b1010101111110100101010111111010010101010110101000010001111001001; end
            14'd7409 : begin out <= 64'b1010101100001001101001010110110110101010100101110010101011001000; end
            14'd7410 : begin out <= 64'b0010011000001010001000101010000010101010010110011010011110011110; end
            14'd7411 : begin out <= 64'b1010011011101100001010010100100110101000100100011010011001110110; end
            14'd7412 : begin out <= 64'b1010100011111101101001101011101110100011100111001010011000001001; end
            14'd7413 : begin out <= 64'b1010010100111101101001101011000000100111000110111010001100100110; end
            14'd7414 : begin out <= 64'b0001111110001011101001011111011000101010101001111010100000000010; end
            14'd7415 : begin out <= 64'b1010000000110010100110101001100110100111010111010001110100010010; end
            14'd7416 : begin out <= 64'b1010010011111001101010010010100110101001001100101010101110101110; end
            14'd7417 : begin out <= 64'b0010011000001100100111011110011110101010001101011010100010110111; end
            14'd7418 : begin out <= 64'b0010100000111010101010111100100000100011101101000001101011010100; end
            14'd7419 : begin out <= 64'b0010010101011011001010001101010110101010111101110010001101101011; end
            14'd7420 : begin out <= 64'b0010101011001011001010011110001110101011111101110010010001110011; end
            14'd7421 : begin out <= 64'b1010101010100000001001100010111110100001110110001010101011111001; end
            14'd7422 : begin out <= 64'b1010101110011001101010100101010110101011110010101010100111111011; end
            14'd7423 : begin out <= 64'b0010010011110001001010100001111110101000101101110010011000110000; end
            14'd7424 : begin out <= 64'b0010100010010000101001000101110010101001100100011010101100000101; end
            14'd7425 : begin out <= 64'b1010011011111110000110001001000000101001111101101001110000011001; end
            14'd7426 : begin out <= 64'b1010100010100000001010100111001010101000100111110010101011010111; end
            14'd7427 : begin out <= 64'b1010010010010111001001101000000010100100110001100010001001010111; end
            14'd7428 : begin out <= 64'b1010010111101100000110000001001110101010100111010010011011011111; end
            14'd7429 : begin out <= 64'b0010100011000111101010101000101010101000110111010010010101101110; end
            14'd7430 : begin out <= 64'b0010100011001101101010101100101000011010001100000010101111000100; end
            14'd7431 : begin out <= 64'b0010100010111000001010111101100110101001010001000010101110000001; end
            14'd7432 : begin out <= 64'b0010010010000000101001111110011110100110100000001010101111001100; end
            14'd7433 : begin out <= 64'b1010100010010111001010010000001010100101110010001010010001110110; end
            14'd7434 : begin out <= 64'b0010101011000001101010111010100010011011011100011000011100100000; end
            14'd7435 : begin out <= 64'b0010100111100110101010000011110010101010000000010010011001000010; end
            14'd7436 : begin out <= 64'b0010100010011001001001100011101010100100100000110010011111000000; end
            14'd7437 : begin out <= 64'b0010011000100101101010001110101110101000011011010010101110101000; end
            14'd7438 : begin out <= 64'b0010011111000000001000101100000010100000000010011010010101011100; end
            14'd7439 : begin out <= 64'b0010010110000110000111100101111110011110110010011010101000110011; end
            14'd7440 : begin out <= 64'b1001100101001000001010111110001100011111010111101001110110110011; end
            14'd7441 : begin out <= 64'b0010100000101000001000011010001000011000110110010010000001011110; end
            14'd7442 : begin out <= 64'b0010100101000101000110000011001100011110011001110010101100001100; end
            14'd7443 : begin out <= 64'b1010100110100110101000110100110000100000001010111010100010110010; end
            14'd7444 : begin out <= 64'b0010000111010010001010001100001010101011101100011010000000010110; end
            14'd7445 : begin out <= 64'b1010100110000000001000011110100110101010001001011010100111110110; end
            14'd7446 : begin out <= 64'b1010100100100010001010100100110000100001001101101010101110101110; end
            14'd7447 : begin out <= 64'b0010100110100100001001110011011010010101011001101010101101111001; end
            14'd7448 : begin out <= 64'b1010010110110101101010111100010000101010101101100001111110000011; end
            14'd7449 : begin out <= 64'b0001100000111010101010110100110000101010001100000010001000100111; end
            14'd7450 : begin out <= 64'b1010101011111100101010100001100000101000100000101001111010111100; end
            14'd7451 : begin out <= 64'b1010010111001010001010010100001100100110000001100010101011100110; end
            14'd7452 : begin out <= 64'b0010100011101110101010111001100110100111110010000010011111110010; end
            14'd7453 : begin out <= 64'b0001011010011000001000111101110000101010100010111010011010101010; end
            14'd7454 : begin out <= 64'b0010100101010011101010101000011000011001010001111010100011111101; end
            14'd7455 : begin out <= 64'b1010100010110110001010001000100000101000111011010010010001110101; end
            14'd7456 : begin out <= 64'b0010010110000100101001101101100100100010110010001010101001010001; end
            14'd7457 : begin out <= 64'b0010100011101101001010010100111100101001001111111010001101011010; end
            14'd7458 : begin out <= 64'b1010100110110011001001110000000100101010110000111010000101100000; end
            14'd7459 : begin out <= 64'b0010011100110011001010101100001000100110011001010010011010001001; end
            14'd7460 : begin out <= 64'b0001111101001011101010101110100000011111000001101010010010111100; end
            14'd7461 : begin out <= 64'b0010101100001111001010110111111110100101110011001010011011000000; end
            14'd7462 : begin out <= 64'b1010010100011101101000011000111010011100011000010001111010011101; end
            14'd7463 : begin out <= 64'b1010100011001011001010110110100110100001100110000001011011010100; end
            14'd7464 : begin out <= 64'b1010011100001110001000101110000010101000101000111010100111101110; end
            14'd7465 : begin out <= 64'b1010100111000000001000100110001010101010111101111001101111101100; end
            14'd7466 : begin out <= 64'b0010100101111011000110101111111100101000101100101010101111001111; end
            14'd7467 : begin out <= 64'b0010101010011100101010110010001010010111110100110010101101011000; end
            14'd7468 : begin out <= 64'b1010001111011011001010011110010000010101101011110001101011001011; end
            14'd7469 : begin out <= 64'b0010000101010111000110110110100110101011111111010010101000101101; end
            14'd7470 : begin out <= 64'b1010010110010011001010010100101110101001110011010010011110010010; end
            14'd7471 : begin out <= 64'b0010011001000100100110011110000110101000000101000010101001101011; end
            14'd7472 : begin out <= 64'b1010100111101001000111001010100110101000111000110010011000100000; end
            14'd7473 : begin out <= 64'b1010011000101101100110001011100000101001111010000001111111100000; end
            14'd7474 : begin out <= 64'b1010101001110011101001010111111000100100011111001010100011011110; end
            14'd7475 : begin out <= 64'b0001011111100100001010101110001100101001111000111010010101111011; end
            14'd7476 : begin out <= 64'b1010101101100110101000100110111000100010110000110010010000001111; end
            14'd7477 : begin out <= 64'b0010011110111110001010000110111100101010101110010010100110011110; end
            14'd7478 : begin out <= 64'b1010010010111001001010111110110100101001101011110010101010110100; end
            14'd7479 : begin out <= 64'b1010101000001010001010101001101000011100101111111010010000010110; end
            14'd7480 : begin out <= 64'b0010000101110000001010001111110100001101000010001010011101100000; end
            14'd7481 : begin out <= 64'b0010100010110010001010010111100110100100100110101010101011110100; end
            14'd7482 : begin out <= 64'b0010011010010000001010010001111110011011011000001010010000011100; end
            14'd7483 : begin out <= 64'b1010101111000100100111110000110100101011000011101010100001111000; end
            14'd7484 : begin out <= 64'b0010101101100111100110010011010110101011011111100010011100011100; end
            14'd7485 : begin out <= 64'b0010010000001100101001011001010110011100001101000010100101101010; end
            14'd7486 : begin out <= 64'b0010100101010111101010110011101010100001100011110010011111010110; end
            14'd7487 : begin out <= 64'b0010100100000100101010100111100110100110010110110001110010000101; end
            14'd7488 : begin out <= 64'b1010100001010110001010010001011000101011001100110010100000110110; end
            14'd7489 : begin out <= 64'b0010110000100000101010010000010110101000011110000010101010001001; end
            14'd7490 : begin out <= 64'b0010010010110000101010010101110000101001101100011001101101010111; end
            14'd7491 : begin out <= 64'b1010011110000001101010000001100000101000100000101001110000010010; end
            14'd7492 : begin out <= 64'b1010100101111101001001000011110000101011101001001010011010100001; end
            14'd7493 : begin out <= 64'b1010010011101101101001110011000000101000001110100010100010111111; end
            14'd7494 : begin out <= 64'b0001111010010100001010100101011100100110010010100010100101010000; end
            14'd7495 : begin out <= 64'b0010100110111101001010100101011000011011010011101010100001001100; end
            14'd7496 : begin out <= 64'b0010100100010101101010111110000000011001101000010010010010010001; end
            14'd7497 : begin out <= 64'b0010101001000100101001000110011010011001000111111001101111010011; end
            14'd7498 : begin out <= 64'b0010001010111101101001101011011100100101101011010010010101111110; end
            14'd7499 : begin out <= 64'b1001100011001000101010100011100000011011100110111010100001011101; end
            14'd7500 : begin out <= 64'b1010101001110010001000100001011110101011111110000010100100110100; end
            14'd7501 : begin out <= 64'b0010100111100111001010100110001010101000000100100010100001101010; end
            14'd7502 : begin out <= 64'b1001110110011100001001001110111010100110111011000010000110011100; end
            14'd7503 : begin out <= 64'b1010100001000000100110010100010110100001111000100010100110100011; end
            14'd7504 : begin out <= 64'b1010010000011101101001011111111100101011001001111001100111000101; end
            14'd7505 : begin out <= 64'b0010001011000101001000011001111010100110000110111010001000110010; end
            14'd7506 : begin out <= 64'b1010101111100101101001101001101010101010100100111010010111101111; end
            14'd7507 : begin out <= 64'b0010100000110110101010010011110100101000010001100010001011100110; end
            14'd7508 : begin out <= 64'b0010100101000110001010100100010100100111001011011010100000010101; end
            14'd7509 : begin out <= 64'b0010101000101011101001011010101000101011100001110010011010100000; end
            14'd7510 : begin out <= 64'b0010010111000110101001001110011000100000001100011010101010001101; end
            14'd7511 : begin out <= 64'b0010101000110011101010010011001000011001001110101010100100000101; end
            14'd7512 : begin out <= 64'b0010100110001001101001110101011000101000001101101010000111001011; end
            14'd7513 : begin out <= 64'b1001110000011100001010010110010100101001010101000010011011000100; end
            14'd7514 : begin out <= 64'b0010101100001010001001011011111110101100001101010010011100011000; end
            14'd7515 : begin out <= 64'b1010011100100000101001000010000010101001111101000010011100010011; end
            14'd7516 : begin out <= 64'b1010100101001001001010101001100010100111011001000010101111000100; end
            14'd7517 : begin out <= 64'b0010101001100000101010010111011100101000101100110010010100000100; end
            14'd7518 : begin out <= 64'b1010101001000100001010010110000110100101000101010010100010111010; end
            14'd7519 : begin out <= 64'b1010100001100010100111010010011110101011000000000010000010001001; end
            14'd7520 : begin out <= 64'b1010001100010101001010010001000110101001001101100010001010101011; end
            14'd7521 : begin out <= 64'b1010000110110101001010100101100000100110110110111001111110100000; end
            14'd7522 : begin out <= 64'b0010010010100110001010011110100110011100010110101010000111011000; end
            14'd7523 : begin out <= 64'b1010000110111001001010100101000010100110000101001010101101011111; end
            14'd7524 : begin out <= 64'b1010101100101100001000011000011010011010110110100010101111011100; end
            14'd7525 : begin out <= 64'b1010100100100110001010001111001000101001110101111010100011111000; end
            14'd7526 : begin out <= 64'b0010101101101101001001110101110110100110010111101010101001001011; end
            14'd7527 : begin out <= 64'b1010101001001001000101011010011100011101111110001010101111100000; end
            14'd7528 : begin out <= 64'b0010000011000011101010101001011010011011011010001010100101110111; end
            14'd7529 : begin out <= 64'b1010100100111010101001110011010000100001010100111010101011001111; end
            14'd7530 : begin out <= 64'b1010000100101001101000101101011110101001101011101010010000111110; end
            14'd7531 : begin out <= 64'b0010101011001101001010101000101110100100000110100010010001100011; end
            14'd7532 : begin out <= 64'b0010101001111010101010011110101110101000100001100010010010000101; end
            14'd7533 : begin out <= 64'b0001111111100110100101000110111110101010000101111001110111000111; end
            14'd7534 : begin out <= 64'b0010100110011001000111001011100010101001110000000010011101010100; end
            14'd7535 : begin out <= 64'b0010100101011000000101000110011110101001101100101010000001101111; end
            14'd7536 : begin out <= 64'b0010001101001100001010110110011010101010001000011010100011010001; end
            14'd7537 : begin out <= 64'b1001110011111000101001100000010010011100000101111010011010001111; end
            14'd7538 : begin out <= 64'b0010000010000111001010000110000010100110110011000010101110110011; end
            14'd7539 : begin out <= 64'b0010011011000001001001100010111000100110110100111010011001010011; end
            14'd7540 : begin out <= 64'b1010101011100001001000001110001110100011011001110010101001100010; end
            14'd7541 : begin out <= 64'b0010100110011000101010010110010110011000100010001010011010000011; end
            14'd7542 : begin out <= 64'b0010101010101110101000100010001010101000000111111010101101101011; end
            14'd7543 : begin out <= 64'b0010100010001100100111000001011100011111111001010010010101000010; end
            14'd7544 : begin out <= 64'b1010000100110011101001000101110100100101011111111010101010100101; end
            14'd7545 : begin out <= 64'b0010101011001000101010000010011010011011111101101010100110001110; end
            14'd7546 : begin out <= 64'b0010101000100010001010000111001000101000000111001010101000000010; end
            14'd7547 : begin out <= 64'b0010011011010000001001001011110100101011100011001010100110101000; end
            14'd7548 : begin out <= 64'b0010101010111000101000000100110100101001010110000010100110100110; end
            14'd7549 : begin out <= 64'b0010101111100000101010000001010110101011000100101010011011110110; end
            14'd7550 : begin out <= 64'b0010100110001001001010101101100110100111110111110001011111110000; end
            14'd7551 : begin out <= 64'b0010101001101111100111100001110010101001111010101010011010010011; end
            14'd7552 : begin out <= 64'b1010010000100101001010011111001100101011111111000010010101000100; end
            14'd7553 : begin out <= 64'b0010001111111011000111110101101100100000011000001010000110000000; end
            14'd7554 : begin out <= 64'b0010100000011101001010001010010010101000111111110001101111111110; end
            14'd7555 : begin out <= 64'b0010000000000100001001011100000110101010110111110010101100001110; end
            14'd7556 : begin out <= 64'b0001101000010010000111010000011000101010111011000010100111101001; end
            14'd7557 : begin out <= 64'b1001111100001011101001010101010000100110110101011010100001111011; end
            14'd7558 : begin out <= 64'b1010011100001111001010010101111000101010011010100010000011001110; end
            14'd7559 : begin out <= 64'b0010100011100000101010001101001010100111000111000001110011110110; end
            14'd7560 : begin out <= 64'b0010011011000111001010100001011010101010111111101010101001000011; end
            14'd7561 : begin out <= 64'b0010100001111011001010111000111010100110111001110010010000111111; end
            14'd7562 : begin out <= 64'b0010011110101011101010101000001000100000101011011010100010001110; end
            14'd7563 : begin out <= 64'b0010101011011111001001001100000110101011101110001010100111001001; end
            14'd7564 : begin out <= 64'b0010100000011100001000001010110110011100110001000001101101111110; end
            14'd7565 : begin out <= 64'b1001111110001111100101001100110100100110101100100010101011100000; end
            14'd7566 : begin out <= 64'b1010101100000000001010100101001110100110111101101001101010000110; end
            14'd7567 : begin out <= 64'b0010101101101000001001000000010000011111100001111010010010100101; end
            14'd7568 : begin out <= 64'b0010100000010100100111110100110100010100111011011010101101010011; end
            14'd7569 : begin out <= 64'b1010001001001100000111001100000000100001110101101010110000010111; end
            14'd7570 : begin out <= 64'b0010010011000110101000001010001110100101000101111001110000111010; end
            14'd7571 : begin out <= 64'b0010101010101111101000010011110110100100011111001010101101111101; end
            14'd7572 : begin out <= 64'b1010100100011110101010111101101000100011010001011010011101000111; end
            14'd7573 : begin out <= 64'b0010010111111100001010010111000000100010111110011010000011000001; end
            14'd7574 : begin out <= 64'b1010011110010111001010011011011110100101110111110010000011010101; end
            14'd7575 : begin out <= 64'b0010001011000111101001100010100110100111011100111010011110000011; end
            14'd7576 : begin out <= 64'b1010100100100111101001100000111100101001111000010010101001101111; end
            14'd7577 : begin out <= 64'b0010110001000010101010010010101100010110000110010010101111111001; end
            14'd7578 : begin out <= 64'b1010010111101111001001100100111000100111110110111010011100111111; end
            14'd7579 : begin out <= 64'b1010011100001111100111110010101010101000101011101010101010010100; end
            14'd7580 : begin out <= 64'b1010011100010011001010000110110100101000111110101010000001110001; end
            14'd7581 : begin out <= 64'b0001011100100101001001001000011100011100111000011010101000000001; end
            14'd7582 : begin out <= 64'b1010100101011000001000010100111100100011101010110010100011100000; end
            14'd7583 : begin out <= 64'b0010100010001111001010000111101110101000011111100010101110000101; end
            14'd7584 : begin out <= 64'b1010000010100001101010000000000000100011110110111010100111100011; end
            14'd7585 : begin out <= 64'b0010101110010110001000011100111100101001011011011010010100111011; end
            14'd7586 : begin out <= 64'b1001101100000101000111110111110110100100101100011010100101000000; end
            14'd7587 : begin out <= 64'b0010100010001011000100010010100100100001111101110010101100100011; end
            14'd7588 : begin out <= 64'b0010100000111011101000001110000100100101011011100010101111001100; end
            14'd7589 : begin out <= 64'b1010100111010100001010011101000010001101101011100010101101001101; end
            14'd7590 : begin out <= 64'b0010100101111000100111111110001000100101100000010010100000100101; end
            14'd7591 : begin out <= 64'b0010100011101000100111011001100010101000110001011010011000110111; end
            14'd7592 : begin out <= 64'b1001111011010110001001100000100010011111111101001010101001001100; end
            14'd7593 : begin out <= 64'b0010101101110111101001100001000010101011001010010001110110010100; end
            14'd7594 : begin out <= 64'b0010011100001110001010010101110100100111100111100010100111111000; end
            14'd7595 : begin out <= 64'b0010101001001111101010000010000100100110100111100010101101100001; end
            14'd7596 : begin out <= 64'b0010100101001101001010100101111110101000111010001010010101010111; end
            14'd7597 : begin out <= 64'b0010001100011111101010011011100000101000010101111010011101111111; end
            14'd7598 : begin out <= 64'b0010010000101010100111000111010100100011111001010010101111011111; end
            14'd7599 : begin out <= 64'b1010001100101000000111110010100000100101101000110010101011010111; end
            14'd7600 : begin out <= 64'b1001110111001001101010101111000010101010010110010010100011000000; end
            14'd7601 : begin out <= 64'b0010101011110110101001111101010010101010110011111010101000101110; end
            14'd7602 : begin out <= 64'b0010100100100110101001110011010110100100110110001010100101111010; end
            14'd7603 : begin out <= 64'b0000111111011111100110001100100000101001001000001010101111100100; end
            14'd7604 : begin out <= 64'b1010100000100000101000010100101100101011000001111010010010000101; end
            14'd7605 : begin out <= 64'b0010101001011111001001100101111000101010110101110010101100001010; end
            14'd7606 : begin out <= 64'b0010101100000111001010010000000100101001111101101010101010100000; end
            14'd7607 : begin out <= 64'b1010101010110011101000000101001010101000010011110010100100001011; end
            14'd7608 : begin out <= 64'b0010001100100000001010110101111010100101001101100010010111100101; end
            14'd7609 : begin out <= 64'b0010100100001100001010001100010010101001001000110001100100110110; end
            14'd7610 : begin out <= 64'b1010001010111001001010111101001010100101101111101010101111101111; end
            14'd7611 : begin out <= 64'b1001101110010011101010001111001000101001000100011010100100011010; end
            14'd7612 : begin out <= 64'b0010001111111011001000111011100000100000000101000010011011011100; end
            14'd7613 : begin out <= 64'b1010010110101101101010111011100110101000001110001001110101011001; end
            14'd7614 : begin out <= 64'b0010101111110110000111000010000010101010110000000010101101010110; end
            14'd7615 : begin out <= 64'b1010011101010100101010000001100010100101100111110001111111111100; end
            14'd7616 : begin out <= 64'b0010001001100011101010111000001110100101110001001010101010010001; end
            14'd7617 : begin out <= 64'b0010001100110011101001001010000010101010110011110010100001111101; end
            14'd7618 : begin out <= 64'b1010011011011110001001000100110100100111000011001010100010111011; end
            14'd7619 : begin out <= 64'b0010000100101111101010100100010010100101001001111010100111011111; end
            14'd7620 : begin out <= 64'b1010101110000001100111010011100100100110001001001010010110000101; end
            14'd7621 : begin out <= 64'b0010101011111111001001100000001010010101111111011010100000011010; end
            14'd7622 : begin out <= 64'b0010011001100011001010111110111000100001000000111010100001110011; end
            14'd7623 : begin out <= 64'b1010100111011011101010000010110000011010100100011010000000000110; end
            14'd7624 : begin out <= 64'b1010011100100111101001000011011110100111000100111010101100011011; end
            14'd7625 : begin out <= 64'b0010100001010010101010110111100000100111010110010010100001001111; end
            14'd7626 : begin out <= 64'b1010100001001100001010001110000100101010011111001010101101010111; end
            14'd7627 : begin out <= 64'b0010100100010000101001110100011100100111011110001010100001110100; end
            14'd7628 : begin out <= 64'b1010011100111011101010011011101100100100001101001010101010011011; end
            14'd7629 : begin out <= 64'b1010101000011001100101101101110110011110001010110001110001001001; end
            14'd7630 : begin out <= 64'b1010100111100011101010101110011010100101001010011010101100101011; end
            14'd7631 : begin out <= 64'b1010101100101001101001100010101010101000101110100010100101010110; end
            14'd7632 : begin out <= 64'b1010101101001011001000011000010100100111011110010010101011110000; end
            14'd7633 : begin out <= 64'b1010000000011110001010000111111100011100110001101010101011011110; end
            14'd7634 : begin out <= 64'b0010101101111110000111100000001000101001100010010001110111001001; end
            14'd7635 : begin out <= 64'b0001110111011001101001100101111110101000000010000010101101100000; end
            14'd7636 : begin out <= 64'b1010010000101100001010010010010010100100100000100001100011110000; end
            14'd7637 : begin out <= 64'b0010101110000100001001010110110010101001111010010010010001110110; end
            14'd7638 : begin out <= 64'b1010101110000100101010110011001010011010111010100010001010011011; end
            14'd7639 : begin out <= 64'b1010011011101100001010010001100100100001100000001010001011110010; end
            14'd7640 : begin out <= 64'b1010101001001011001010011111011000101011100100000010100100001011; end
            14'd7641 : begin out <= 64'b0010100110001001001010000100001010101000111001011001100110101100; end
            14'd7642 : begin out <= 64'b1010001000111110101001001100111010100000110100010010001001011000; end
            14'd7643 : begin out <= 64'b1010001110100100101010110010011110101010000110011010101010100101; end
            14'd7644 : begin out <= 64'b1010011111111010100110111011001110100011010110000001001110001010; end
            14'd7645 : begin out <= 64'b0010101111111010001001110110111000100111110100010010100101001111; end
            14'd7646 : begin out <= 64'b0010101010001000100101111101101100100001010111011010100101000011; end
            14'd7647 : begin out <= 64'b0010100110010011001000100101001000101010100001101010011010100111; end
            14'd7648 : begin out <= 64'b1010011010000110001010001110011110100010100001000010011100100000; end
            14'd7649 : begin out <= 64'b1010010101110001000111000001110000101001001011011010101000000101; end
            14'd7650 : begin out <= 64'b0010011001010111001010011001001100101000001011011010100101000100; end
            14'd7651 : begin out <= 64'b0010011001010111101010100011011000101010100011100001111111110010; end
            14'd7652 : begin out <= 64'b1010010011100111001010100100000000010100010000100010000010010101; end
            14'd7653 : begin out <= 64'b0010001110111000001010000011001010100110010001000010100111010011; end
            14'd7654 : begin out <= 64'b0010000010011010101000100111011010101011000110001010100111110011; end
            14'd7655 : begin out <= 64'b1010011100001011101010111110000010011111110010000010100100100011; end
            14'd7656 : begin out <= 64'b0010011101011110101001001000100000101010101111011010100110110000; end
            14'd7657 : begin out <= 64'b1010101101110111101000011011011000101011001000100010101000101100; end
            14'd7658 : begin out <= 64'b0010101101010010001000110011101010101001100110010010010000010000; end
            14'd7659 : begin out <= 64'b1010100100001100001001101010001000011100110010100010101101010101; end
            14'd7660 : begin out <= 64'b1001100011010110001010101000001000101100000011000001110110101001; end
            14'd7661 : begin out <= 64'b0010101101100110001001010011110110011101011000000001001000000001; end
            14'd7662 : begin out <= 64'b0010100011011110101010101111001100100001001111100010001111000101; end
            14'd7663 : begin out <= 64'b1010100001110101000111101011111100010000110101101010101011100010; end
            14'd7664 : begin out <= 64'b0010010111110000100011000110100000100111101010111010100110011011; end
            14'd7665 : begin out <= 64'b0010011011111111101010100000101110100000000110011010010000100101; end
            14'd7666 : begin out <= 64'b0010010111010110101001001110101000101000101011110010101001011010; end
            14'd7667 : begin out <= 64'b1010100100110111001001010110111110011000101010000010010111010000; end
            14'd7668 : begin out <= 64'b1001110110001100001010100011110010101011111010010010101101101001; end
            14'd7669 : begin out <= 64'b0001111011010100100011010100101000100101001110000001101000101110; end
            14'd7670 : begin out <= 64'b1010000011011111000111011111101110010101000100100010000101000000; end
            14'd7671 : begin out <= 64'b1010011111010001101001101111001010100101010110111010100100101001; end
            14'd7672 : begin out <= 64'b1010011111111000001000000110010000010010110111011010010001101001; end
            14'd7673 : begin out <= 64'b0010011110111111001001111010000000100011111001100010110000001110; end
            14'd7674 : begin out <= 64'b1010101110100011101010010001000100100100110110010010001001011111; end
            14'd7675 : begin out <= 64'b1010100000101010001010001101000010101010110001000001110010100011; end
            14'd7676 : begin out <= 64'b0010100011000010000111011011101110101011110011011010011000110010; end
            14'd7677 : begin out <= 64'b1010011110111001101000110100000000100111100010110010101101101000; end
            14'd7678 : begin out <= 64'b1010100000100110001000000110000110100001110001011010001100110001; end
            14'd7679 : begin out <= 64'b1010101100111101001001011110000000101100001010011010100111010110; end
            14'd7680 : begin out <= 64'b0010010111011100001001001010111010101010100111111010010101101011; end
            14'd7681 : begin out <= 64'b0010011010111110101001101100011000100010010110101010100001101111; end
            14'd7682 : begin out <= 64'b0010010100001011101010001101011100100100111010100010011100011000; end
            14'd7683 : begin out <= 64'b1010101010101011101010100100111100011101101110000010100011100100; end
            14'd7684 : begin out <= 64'b0010010110110011001000011000011000100011011010011010011001100011; end
            14'd7685 : begin out <= 64'b0010001110001011101001011001010100101011100010110010101000111101; end
            14'd7686 : begin out <= 64'b0010101001100000001010010111100110101000110110101010100101101110; end
            14'd7687 : begin out <= 64'b0010100001100001000110011001111010100010010111111010101001010010; end
            14'd7688 : begin out <= 64'b1010011010101010100100010010111110011101000100111010011000100011; end
            14'd7689 : begin out <= 64'b0010001100101000101010100000000000100100101001101001110101111110; end
            14'd7690 : begin out <= 64'b0010101101001001001001001000001110101011101101111010011101100110; end
            14'd7691 : begin out <= 64'b0001100011010000101010011001101010101001101010110010101111101100; end
            14'd7692 : begin out <= 64'b0010101110011111001010111000001010100110001100110010101000001110; end
            14'd7693 : begin out <= 64'b0010100001110001100111100111000110101000001100001010011110111011; end
            14'd7694 : begin out <= 64'b1010101101010110000111110010110000100100000001000001011000110010; end
            14'd7695 : begin out <= 64'b0010011001110100101001110011000110100110001100110010101010100011; end
            14'd7696 : begin out <= 64'b1010101100011110000110000000100100101001010111101010001110110101; end
            14'd7697 : begin out <= 64'b0010100000001011100111010010011010010011100100100010100010111111; end
            14'd7698 : begin out <= 64'b0010011010100111000111000010001010101001100001110010100111011101; end
            14'd7699 : begin out <= 64'b1001110001111010101010001011011100100010110010011010101000010000; end
            14'd7700 : begin out <= 64'b0010101111100001101001001111000100101000110000111010011001110011; end
            14'd7701 : begin out <= 64'b1001111000010101001001010111010110101000011100101001110101110001; end
            14'd7702 : begin out <= 64'b0010101000100111101010100001111100100101100001111010100111001111; end
            14'd7703 : begin out <= 64'b0010011111101001001001011011011100101000110101011010101111110011; end
            14'd7704 : begin out <= 64'b1010100101110100001010101001001000101000000101100010011100110101; end
            14'd7705 : begin out <= 64'b1010011010000111101001011011011010101011000101010001111011000101; end
            14'd7706 : begin out <= 64'b1010100010101111001010001110100110101000010111101010100010110111; end
            14'd7707 : begin out <= 64'b1010100100000011001010000100111110101011011011101010101000011111; end
            14'd7708 : begin out <= 64'b1010101111111110101010010110001110100100100110111010010010010001; end
            14'd7709 : begin out <= 64'b0010101101001111101000001110000000101001111010111010101000101001; end
            14'd7710 : begin out <= 64'b1010100000010111100011110010100100100101100001111010101001110000; end
            14'd7711 : begin out <= 64'b1001111001000010001010001001111010100101010010110010000101101000; end
            14'd7712 : begin out <= 64'b1010100100001001101010100100001100100111100010110010100100000100; end
            14'd7713 : begin out <= 64'b0010100100010110000111110011010110101010100011001001111000101011; end
            14'd7714 : begin out <= 64'b0010101101111010001010101001011110101001010001001010010101011011; end
            14'd7715 : begin out <= 64'b0010011001111000101010011111110110101001110110100010100001110101; end
            14'd7716 : begin out <= 64'b0001111001111111001001010001001110100111111010010010100101010111; end
            14'd7717 : begin out <= 64'b1010001010000011101010011001110110101000011110110010000000011011; end
            14'd7718 : begin out <= 64'b0010101100101011001010001111010000101001001000100010011111000110; end
            14'd7719 : begin out <= 64'b1010010100111100100111000000000110101011111001000010000010111000; end
            14'd7720 : begin out <= 64'b1010000100111010001010001111100100100100011111010010101110000100; end
            14'd7721 : begin out <= 64'b1010100000011100101010011101001100101001011011010010101000011101; end
            14'd7722 : begin out <= 64'b1010101011101000001010001100000010101001011011001010011110000110; end
            14'd7723 : begin out <= 64'b0010101110011111100111110011010010100010101010110001111000110100; end
            14'd7724 : begin out <= 64'b1010100000101000000111001101100110100110111001010001110010000100; end
            14'd7725 : begin out <= 64'b0010101011101101101001110011111100101010001101100010011100100100; end
            14'd7726 : begin out <= 64'b0010011000101101101010010001100000100010110011110010011111101100; end
            14'd7727 : begin out <= 64'b0010101100101101001010011000111100101011111000001001101010011010; end
            14'd7728 : begin out <= 64'b1010001101100010101000110000100100101000011110000010000011001101; end
            14'd7729 : begin out <= 64'b0001110111001110000110011111011000101011100111011010100110110111; end
            14'd7730 : begin out <= 64'b1010011101100000100110000110110000101000010001101010101000011000; end
            14'd7731 : begin out <= 64'b0010101100111110101010101110101110100001110010001010101111101011; end
            14'd7732 : begin out <= 64'b1010100001001010101001000011011100101011010100000010101000101010; end
            14'd7733 : begin out <= 64'b0010100010001010101010011001000010010111001101100010001110101111; end
            14'd7734 : begin out <= 64'b0001111111101000100110110000010110101010011011100010101100001100; end
            14'd7735 : begin out <= 64'b1010100100100010101001011011111000101001111111010010010001100010; end
            14'd7736 : begin out <= 64'b0010101111101001101010010100100000100011101000100010011110101010; end
            14'd7737 : begin out <= 64'b0010010010001010101010100001101010100110110100101010101100101100; end
            14'd7738 : begin out <= 64'b1010100101101001101010101101110110011001010101000001011110010001; end
            14'd7739 : begin out <= 64'b0010001000101111101010110001110000100010100111011010100100101001; end
            14'd7740 : begin out <= 64'b1010011100001011001010100111011010101010001101110010100110101011; end
            14'd7741 : begin out <= 64'b0001001000001010101001110010111100011101101011000010000010000001; end
            14'd7742 : begin out <= 64'b1010101100100111101010101101101010101000011110011010100100001111; end
            14'd7743 : begin out <= 64'b0010100110010100101001100101010010101000101101100010101000100000; end
            14'd7744 : begin out <= 64'b1010101001101010101010100100010100101010100101100010011001110100; end
            14'd7745 : begin out <= 64'b1001110100011010001010011101010100100011001100000010101010101110; end
            14'd7746 : begin out <= 64'b1010101010100010001010101101110110100010111000101010000011101101; end
            14'd7747 : begin out <= 64'b0001011010100111100111011110010000101010011001011010101000011011; end
            14'd7748 : begin out <= 64'b1010011110001000101010000101011000100000111000100010101000100010; end
            14'd7749 : begin out <= 64'b0010100111010111001010001010110010101000011001000010101000110110; end
            14'd7750 : begin out <= 64'b0001110001101100101010011101001110101100000001101010101101110101; end
            14'd7751 : begin out <= 64'b0010011000001111001001000011111100101001101111011010100111101000; end
            14'd7752 : begin out <= 64'b1010101000010011101010010011001010101000101001011010000101110100; end
            14'd7753 : begin out <= 64'b1010101001101011001010000001111010101001111001111010101000000111; end
            14'd7754 : begin out <= 64'b0010011101001101101011000100011100101000000011001010101110010011; end
            14'd7755 : begin out <= 64'b0010101010000000101010111001100100101011101110011010011001000001; end
            14'd7756 : begin out <= 64'b1010101111001000101001011000000000011110011000101010011111010011; end
            14'd7757 : begin out <= 64'b1010001011100000000111010111010110101001111010001010100111001001; end
            14'd7758 : begin out <= 64'b1010101111000100101000111001000110100010101011100010100110000011; end
            14'd7759 : begin out <= 64'b1010100110010101101010101111110110011100110001010010100000000111; end
            14'd7760 : begin out <= 64'b0010010000100001001001100100100000101001010000010010000110110010; end
            14'd7761 : begin out <= 64'b1010101111110110101010100101001000101011010001000010010110001001; end
            14'd7762 : begin out <= 64'b0001111111011000101001111010010000101011010110011010101110001010; end
            14'd7763 : begin out <= 64'b0010010011000000101010111000001010101001110000101010101111000011; end
            14'd7764 : begin out <= 64'b0010101011010111101001101010011110101011011101101001000110010010; end
            14'd7765 : begin out <= 64'b0010100011011110101000000000010100101000000010111010001101010110; end
            14'd7766 : begin out <= 64'b1010101101011110000111010011010010101000100100111010100111001100; end
            14'd7767 : begin out <= 64'b1010010110100011001010101000100100011110011010001010101010111111; end
            14'd7768 : begin out <= 64'b0010100101010011101010110001011110100100101111011010010000111000; end
            14'd7769 : begin out <= 64'b1010001011101010000111100111001010101000010111010010001100100100; end
            14'd7770 : begin out <= 64'b1010010000010000101010001010100010100001001011000010010011001011; end
            14'd7771 : begin out <= 64'b0010011011001100001010011010001100101011001001101010010001100111; end
            14'd7772 : begin out <= 64'b1010010111111010101010011111010010100110000011110010001001000010; end
            14'd7773 : begin out <= 64'b1010011011010110101000110010011000100001110100111001110110001001; end
            14'd7774 : begin out <= 64'b0010010101010001001000111011100010100010111110000010010111001111; end
            14'd7775 : begin out <= 64'b0010100010110000001010101101101010100111110100010010100000110001; end
            14'd7776 : begin out <= 64'b0010101011010111101001000001110100101010110010101010011001000001; end
            14'd7777 : begin out <= 64'b1001010100101101001010101010101100011101101100010001001010110111; end
            14'd7778 : begin out <= 64'b1010100001010110001000000000010110100110100000111010100100010011; end
            14'd7779 : begin out <= 64'b0010100011110100001000111010001110101011000000011010100110110100; end
            14'd7780 : begin out <= 64'b1001101011110001101010111100001110101000111011000010101100010100; end
            14'd7781 : begin out <= 64'b1010100100110010001010010011110000101011101011110010001011110100; end
            14'd7782 : begin out <= 64'b1010101111111111001010101001110100100111101011111010001000011101; end
            14'd7783 : begin out <= 64'b0010011000100110001010101010100100101010011000111000111110100101; end
            14'd7784 : begin out <= 64'b0010011000001001001010110001001110101011000010000010100110011000; end
            14'd7785 : begin out <= 64'b0010010110011100101001111011001000101011110010100010011110101001; end
            14'd7786 : begin out <= 64'b0010100000110101001010000000101110100110111000111001101100011010; end
            14'd7787 : begin out <= 64'b1010010100110101101001010000010110101001111000010010011100011001; end
            14'd7788 : begin out <= 64'b1010011100101100100111110000010010010101111111010010010010001001; end
            14'd7789 : begin out <= 64'b1010011010011111001001100000011010101010100110101010011000111011; end
            14'd7790 : begin out <= 64'b1010010010000110000111001111110100100100001001111010101111111001; end
            14'd7791 : begin out <= 64'b0010001101110100001001110000011000101011000001011001110001000001; end
            14'd7792 : begin out <= 64'b1010101101010010100110101010000100101000001010111001100010101000; end
            14'd7793 : begin out <= 64'b1001001111000111101010001101101010101001011011101010100101011110; end
            14'd7794 : begin out <= 64'b0010101100010110001001011111111010100101100001011010100111101011; end
            14'd7795 : begin out <= 64'b0001110110001111001001010001001100011100100100100010000001111000; end
            14'd7796 : begin out <= 64'b0010101001001100001000000001110100011110111011011010010001101101; end
            14'd7797 : begin out <= 64'b0010001001000000001010001001110100101000001111000010000100010101; end
            14'd7798 : begin out <= 64'b1010100101011111001010101111001110101000011001000010100010100100; end
            14'd7799 : begin out <= 64'b1010001011011011001010111000011110011010100100001010011110000100; end
            14'd7800 : begin out <= 64'b1010011010101010001010111100000000101001110000010001010110000011; end
            14'd7801 : begin out <= 64'b0010011101001110101010011111000100101001010000110001101000101100; end
            14'd7802 : begin out <= 64'b0010000110100010101011000101000000101001001010111010001100000010; end
            14'd7803 : begin out <= 64'b1010100011111010101010010100101010101011011111011010011010010101; end
            14'd7804 : begin out <= 64'b0010000100010111101001101011010010100101001101110010101010110010; end
            14'd7805 : begin out <= 64'b1010101101111000001001011101111100101011011010011010011100101010; end
            14'd7806 : begin out <= 64'b0010100110111100101001111100100100101011000001011010100101001101; end
            14'd7807 : begin out <= 64'b0010101100010101000001100111011100101011011011001010010100010100; end
            14'd7808 : begin out <= 64'b1001011110000111101010011010001000100100011010011010010011111001; end
            14'd7809 : begin out <= 64'b0010101011111010001000011110101100101011001101100010010111110010; end
            14'd7810 : begin out <= 64'b0010101110110000001010110001100000101011011001011010101000100100; end
            14'd7811 : begin out <= 64'b0010100010100111001010101111011010101011000110011010101000001101; end
            14'd7812 : begin out <= 64'b0010100000000110101001100101101000101010010010011001111010011001; end
            14'd7813 : begin out <= 64'b0010100111000101101010100110001100011111110110111010100000000110; end
            14'd7814 : begin out <= 64'b0010101111011001001010101111101000101010000110000010001100011001; end
            14'd7815 : begin out <= 64'b1010100100100110101010000010001100101010000101110010011000010001; end
            14'd7816 : begin out <= 64'b1010100101001010001001111101101000100100101110100010101000110111; end
            14'd7817 : begin out <= 64'b0010100101100011101010011101110100101010111110110010100110011111; end
            14'd7818 : begin out <= 64'b0010011111101001101010011011101010100111000101000010010011101100; end
            14'd7819 : begin out <= 64'b1010011111001011101010101111001010100010000111000010010110011110; end
            14'd7820 : begin out <= 64'b0010011000001010001000000101011100101011110100111010100100011011; end
            14'd7821 : begin out <= 64'b0010100111001010001010100101010010101001101000101010010000111010; end
            14'd7822 : begin out <= 64'b0010101010001001101000000001111000100101000100111010001101011100; end
            14'd7823 : begin out <= 64'b0010010010000011000111001010000100011100110100101010100101101001; end
            14'd7824 : begin out <= 64'b0010101101000001101010101011000000101001010010111010100101000111; end
            14'd7825 : begin out <= 64'b0010101011100101101010010101101100101010010111010010001010000111; end
            14'd7826 : begin out <= 64'b0010011000010000001010110000010100100101110111111010100110110011; end
            14'd7827 : begin out <= 64'b0010100100000100101010010011011010101001110000000010100010110000; end
            14'd7828 : begin out <= 64'b1010001100111000001000001100101010100011110010111010101000001110; end
            14'd7829 : begin out <= 64'b0010101011100001001001100110110100100101000111100010101110100001; end
            14'd7830 : begin out <= 64'b0010101000000101001010011101100110101000111010111010100011100111; end
            14'd7831 : begin out <= 64'b0010100001010111101010110111011010101011100100001010100000011011; end
            14'd7832 : begin out <= 64'b0010000000000110001001010101110010101001110010111010100010000100; end
            14'd7833 : begin out <= 64'b0010100011001001101010010000101110101000000000000010101110110100; end
            14'd7834 : begin out <= 64'b0010011000010010001001010001001110101010111011011010100000011111; end
            14'd7835 : begin out <= 64'b1010101001111011101001001100100010101010000101100010010010111110; end
            14'd7836 : begin out <= 64'b1010011001101100001001100110101100101000101100100010101100011111; end
            14'd7837 : begin out <= 64'b0010101101110011001010110110100110101000011111011010011100101011; end
            14'd7838 : begin out <= 64'b1010101111110110101001000111000000100110100010100010100011000101; end
            14'd7839 : begin out <= 64'b1010000110001110100111110011101010011110100001000010101001110011; end
            14'd7840 : begin out <= 64'b0010100110110101101010100011111010100010000011011010000001101110; end
            14'd7841 : begin out <= 64'b1010101001101110101010101101111100101010111010001010011110000011; end
            14'd7842 : begin out <= 64'b0010000101111101101000001101110000101010001101010010011000000101; end
            14'd7843 : begin out <= 64'b0001110010011000101001100001011010100101011100110001110101010110; end
            14'd7844 : begin out <= 64'b1010011001011011101010111100100010101011001011100010100101100111; end
            14'd7845 : begin out <= 64'b0010101011011110001011000000111000100110100100100010100111110010; end
            14'd7846 : begin out <= 64'b1010100001101101101001101101101000100100110001010010100110111010; end
            14'd7847 : begin out <= 64'b0010101110001001001010001101100110101001111100110010010111011011; end
            14'd7848 : begin out <= 64'b0010100000111001001000001010011110100011010011010010011001001110; end
            14'd7849 : begin out <= 64'b1010100111110000001010010101110010101010100001011010101110100011; end
            14'd7850 : begin out <= 64'b0010001000000010001001011111000110100101111101010010100001100101; end
            14'd7851 : begin out <= 64'b0010100001100110000111110101000000011101100000110010101001001111; end
            14'd7852 : begin out <= 64'b1010101100100110001001010000000100101000111000100010101011011111; end
            14'd7853 : begin out <= 64'b0010101001011111101010011110100010100111011001100010101111011110; end
            14'd7854 : begin out <= 64'b1010101100011101001010111111011010101000011101111010011000011100; end
            14'd7855 : begin out <= 64'b1001111000000001101010111001011000101010011110001010100111111001; end
            14'd7856 : begin out <= 64'b1010010010111000101010001111101110101001010001110010010101011110; end
            14'd7857 : begin out <= 64'b0010101101101011000111110010000010101011110000001010010010110010; end
            14'd7858 : begin out <= 64'b0010001110011101001001011110111110011100111000110010100001001111; end
            14'd7859 : begin out <= 64'b0010101010110000101001001011100100100110110011101010101011000111; end
            14'd7860 : begin out <= 64'b0010101011010010001001011110000000011111001011110010100101000100; end
            14'd7861 : begin out <= 64'b0010010110001001101010111011111100010000111100100010101011010111; end
            14'd7862 : begin out <= 64'b1010010100011000101001011100000100101001011100000001111101011001; end
            14'd7863 : begin out <= 64'b1010100100101010100111111101000110101000111001100010011001001001; end
            14'd7864 : begin out <= 64'b1010101100110110101010010101011000100001110010010010011000011111; end
            14'd7865 : begin out <= 64'b0010100011101101101000001000100010101011010111001010011011100010; end
            14'd7866 : begin out <= 64'b0010011011010100101001001001000100101011110011010001100000001001; end
            14'd7867 : begin out <= 64'b0010100000110111001000001101100000101000101101101010100100101010; end
            14'd7868 : begin out <= 64'b1010100001011011100101101101111010101010101001111010011001010001; end
            14'd7869 : begin out <= 64'b1010100111100111101010101000110110100100110100001010100001110000; end
            14'd7870 : begin out <= 64'b1010101010010110001010011110010100101011111111011010011111110101; end
            14'd7871 : begin out <= 64'b1010100101010110101010111101011100100000010110011010101110000001; end
            14'd7872 : begin out <= 64'b0010100010011111001010001010101010101010110011000010000110001010; end
            14'd7873 : begin out <= 64'b1001111110111011101010010001110110101000110101000010101000111110; end
            14'd7874 : begin out <= 64'b1010010000010111101001000110100010101011111000001010100001110010; end
            14'd7875 : begin out <= 64'b0010000010110110101011000000010010100100010101011010010001001110; end
            14'd7876 : begin out <= 64'b0010011010101010101000000101101000100011100010101010000000001100; end
            14'd7877 : begin out <= 64'b0010100000111100101001101110010110101011100110011010100101100111; end
            14'd7878 : begin out <= 64'b0010011001101110101010111100111010010111100001000010101010110001; end
            14'd7879 : begin out <= 64'b0010000010011000001000111001101000101011001001011010100011100110; end
            14'd7880 : begin out <= 64'b0010101111111100101001000101000110100001010101001010100001100000; end
            14'd7881 : begin out <= 64'b1010100110110001001001110100110000101011001111101010010111111000; end
            14'd7882 : begin out <= 64'b1010100100000010000111011111010100101001110000111001100110100011; end
            14'd7883 : begin out <= 64'b0010101001000001001010111101010110101011010001110010000001000110; end
            14'd7884 : begin out <= 64'b0010100011010111001010011010011010011111010111010010100011101111; end
            14'd7885 : begin out <= 64'b1010010101011000101001000101001110101010011010000010100010101100; end
            14'd7886 : begin out <= 64'b1010100000110011101000011001101010100111100001001010001101111111; end
            14'd7887 : begin out <= 64'b1010100101110111001010100010110010011110010100011010101110010100; end
            14'd7888 : begin out <= 64'b1010100101111001101010101001101110100111011010101010101100010011; end
            14'd7889 : begin out <= 64'b0010101011000100001010101100101000101010110111000010101000000101; end
            14'd7890 : begin out <= 64'b0001010101111011101010000100001110101001110100011010101111000011; end
            14'd7891 : begin out <= 64'b0010100111110110001010011010001110101010101001100010101000111000; end
            14'd7892 : begin out <= 64'b1010100011110000001010110001101100011011100100100010100100100000; end
            14'd7893 : begin out <= 64'b0010101011000001001011000000101010101011010100001010001110011101; end
            14'd7894 : begin out <= 64'b0010010101011101101010001010001010011111110111111010010010000100; end
            14'd7895 : begin out <= 64'b1010101110000101101010110001000000101010011101011010010111000011; end
            14'd7896 : begin out <= 64'b0010100001010110101010101010011000101010001100010010001001001110; end
            14'd7897 : begin out <= 64'b0010101000110101101010011100101100101010111110001010010010001010; end
            14'd7898 : begin out <= 64'b0010000101010001101010011110011100011000111110010010101011001111; end
            14'd7899 : begin out <= 64'b1010010001000110001001010111000100100101101111111010001100010100; end
            14'd7900 : begin out <= 64'b0010011111101111000111000010101010100111110110011010011011110000; end
            14'd7901 : begin out <= 64'b0001101100010010000111010000011000100101111101101010101001110111; end
            14'd7902 : begin out <= 64'b0001111101111001101001001000010010101010001111000010011001001101; end
            14'd7903 : begin out <= 64'b1010101111111010100111110000010100010110111000011010011000010001; end
            14'd7904 : begin out <= 64'b0010100101011101101010100100010000101001110010011010011101100101; end
            14'd7905 : begin out <= 64'b1010100101001001001000010110011110100101111100111010010101011110; end
            14'd7906 : begin out <= 64'b1010101011011110101010001111110100101011010100010010011011001001; end
            14'd7907 : begin out <= 64'b1010100000110000001001000101110100100111101011011010101000100111; end
            14'd7908 : begin out <= 64'b0010010011110001101010000001100110101000000011011010100110000001; end
            14'd7909 : begin out <= 64'b1001110111010011101001101111001100101000101110100010101000000111; end
            14'd7910 : begin out <= 64'b1010100010100001101010000110101100011111101100101010101111110111; end
            14'd7911 : begin out <= 64'b1010100111111110001001100011111110101000000101100010000000000001; end
            14'd7912 : begin out <= 64'b1001111110011111101010101011100110010110111111001010100100000011; end
            14'd7913 : begin out <= 64'b0010100000101111001001100101011110010000010111000010000011011110; end
            14'd7914 : begin out <= 64'b1010100100111101101010100101010010100101011000111010010011100001; end
            14'd7915 : begin out <= 64'b1010101100100001001001001101111110100010110100011010101100111000; end
            14'd7916 : begin out <= 64'b1001110010010001001010110011011010101010101010111010010101110011; end
            14'd7917 : begin out <= 64'b0010100111011011001010100111111000010111110011001010100111110110; end
            14'd7918 : begin out <= 64'b1010100010101111101000010001101010100001001111010010101001011010; end
            14'd7919 : begin out <= 64'b0010011100100001001001100000000110101011010010001001100111010001; end
            14'd7920 : begin out <= 64'b1010011100000000101000010101110000100001111000000010001101010101; end
            14'd7921 : begin out <= 64'b1010101110010100101001110001111000101011111110110001111010110100; end
            14'd7922 : begin out <= 64'b0010001000001110100111110000001110101000110000001010000111000100; end
            14'd7923 : begin out <= 64'b1010101100101010101001000001010000101001001100111001110101001001; end
            14'd7924 : begin out <= 64'b1010011011111010101010010001110100100001111111101010100111001010; end
            14'd7925 : begin out <= 64'b1001101101010111001001010000110000101001100111110010101100011111; end
            14'd7926 : begin out <= 64'b1010101110100110101011000100011110101000100011010010001000010010; end
            14'd7927 : begin out <= 64'b0010011000011100101001010000010100100111010111101010001010001101; end
            14'd7928 : begin out <= 64'b1010101000010001001010100010111100100000010011110010000110010011; end
            14'd7929 : begin out <= 64'b0010010110010101000111001111101000101000100010011010100111100010; end
            14'd7930 : begin out <= 64'b0001100011110101101001110010010110101000111101100010101101000101; end
            14'd7931 : begin out <= 64'b1010100001100111001010101010110100101010100110011001111000001011; end
            14'd7932 : begin out <= 64'b0010011001111011101010101010101110101001011111111010011101000100; end
            14'd7933 : begin out <= 64'b0010010101000011101010001001100010101001101011101010100011001111; end
            14'd7934 : begin out <= 64'b0010101000010011001010010101110110100000111110110010010110111011; end
            14'd7935 : begin out <= 64'b0010101100101110100111011000101110011110111001001010100101010000; end
            14'd7936 : begin out <= 64'b1010011101101011001010001101100000100110011010101010100001010100; end
            14'd7937 : begin out <= 64'b0001000000001101101010110001011100100100111001100010101001011100; end
            14'd7938 : begin out <= 64'b1010101110000011001000111110001100100110010001111010101111110101; end
            14'd7939 : begin out <= 64'b0010010011001100100111011110101000010100100001100010110001011110; end
            14'd7940 : begin out <= 64'b1010100000001010101001101010010010101001010110101001001001100010; end
            14'd7941 : begin out <= 64'b1010011010110110100111011101011010101011100010010001001111111110; end
            14'd7942 : begin out <= 64'b1001110101000001101010010001000000010111010110110010100101111000; end
            14'd7943 : begin out <= 64'b0010010110101101001010000010110000101001111100011010100000001100; end
            14'd7944 : begin out <= 64'b1001110110010000001010010011000100100110101110101010101011000001; end
            14'd7945 : begin out <= 64'b0010001000011011101000110001110110100111110100100010100110111110; end
            14'd7946 : begin out <= 64'b0010100000100010001010110111000000100100110100000010110000010111; end
            14'd7947 : begin out <= 64'b1010011001101101101010101000100000101000011011110010101001001001; end
            14'd7948 : begin out <= 64'b0010100001000011101010000101000010101001000101100001100100011011; end
            14'd7949 : begin out <= 64'b0010100101110110001010111110101110101010010001001010101011101101; end
            14'd7950 : begin out <= 64'b0010101010001011101001010110001000101010111011011010101000100000; end
            14'd7951 : begin out <= 64'b1010010101010101101000100010010110101010010000010001000011001110; end
            14'd7952 : begin out <= 64'b1010000101001011001000000010101100101010111010011001110100110010; end
            14'd7953 : begin out <= 64'b1010101111000111101010110101111100100111000010110010010101000000; end
            14'd7954 : begin out <= 64'b0010100001011010101010011010101110101010010000001010101011000010; end
            14'd7955 : begin out <= 64'b0010100000111110001010110011001010101000000101001010101000010011; end
            14'd7956 : begin out <= 64'b0010000101001001000100111011110000101001100011111010001010110100; end
            14'd7957 : begin out <= 64'b1010101110111111101010000110011010101001010110100010100001001101; end
            14'd7958 : begin out <= 64'b1010100000001110000111111110101110101010111101110010011001010000; end
            14'd7959 : begin out <= 64'b1010101001010001101010001100000110101001011010111010101101100111; end
            14'd7960 : begin out <= 64'b1010101100000110101010110101001100100000010011011010100000111001; end
            14'd7961 : begin out <= 64'b0010100101010101001010001010010110101001000000100010011111110000; end
            14'd7962 : begin out <= 64'b1010011110100000001001011000111110100101101000100010101000001100; end
            14'd7963 : begin out <= 64'b0010100000100111101010111110000110100101000001010010101001100011; end
            14'd7964 : begin out <= 64'b0010000011101000001000001000011110100011011101110010010010011000; end
            14'd7965 : begin out <= 64'b0010110000001011001000001101110100101001100111101010000111000100; end
            14'd7966 : begin out <= 64'b0010100001010100001001100110011010101001101100010001101110000101; end
            14'd7967 : begin out <= 64'b0010001000101110101010100100111110100110011010011010011101110101; end
            14'd7968 : begin out <= 64'b1010000010111011101010001010101000100111111001010001011000010001; end
            14'd7969 : begin out <= 64'b0010101001111001001010100010110100101011010001101010010000011001; end
            14'd7970 : begin out <= 64'b1010100000001010101010011011010110101010100101011001111111101100; end
            14'd7971 : begin out <= 64'b0010100110001100101010000011000100101000101110001010010100100001; end
            14'd7972 : begin out <= 64'b0010100001011110001010011111110000101011001011110001111101001100; end
            14'd7973 : begin out <= 64'b1010101011110001001000100111101110101010100101100010101011110000; end
            14'd7974 : begin out <= 64'b0010100101001110001000101011110000101010111001010010011001100000; end
            14'd7975 : begin out <= 64'b0010011110100110001010010100010010101000111011010010000110001111; end
            14'd7976 : begin out <= 64'b0010101100011110101010111110010100010100000001110010011101010011; end
            14'd7977 : begin out <= 64'b1010000111100001001010100111001010101011101100000010001000011011; end
            14'd7978 : begin out <= 64'b1010001100000010001001100111000110101011101100110010000111111111; end
            14'd7979 : begin out <= 64'b1010010100110100101001101011101010100000111010010010100101111010; end
            14'd7980 : begin out <= 64'b0010000011011101001010111001111110100110111110010010100110110001; end
            14'd7981 : begin out <= 64'b0010001111111011100100110001011000100000101011100010101001110100; end
            14'd7982 : begin out <= 64'b1010101110110011101001101000000100011110110010011010000100010100; end
            14'd7983 : begin out <= 64'b0010011011011010001010010010011000011001010101001010100000011101; end
            14'd7984 : begin out <= 64'b1001111000001100101010100111011000101010011001101001111001100100; end
            14'd7985 : begin out <= 64'b0010101010101110101001010011101000101000000000011010101100010101; end
            14'd7986 : begin out <= 64'b0010100011000100101010000100010010011110100010000010101000011111; end
            14'd7987 : begin out <= 64'b1010100110001100001010110000010000101001100000100010010110111100; end
            14'd7988 : begin out <= 64'b1010100001010101001010110111100100010110110101011010000011010010; end
            14'd7989 : begin out <= 64'b1010100111011010001010111111100000101001110110101010100011111100; end
            14'd7990 : begin out <= 64'b0010100010010101001001100100001110100111011000001010011000100110; end
            14'd7991 : begin out <= 64'b1010101000010000101000100011101010101000011001011010011100110001; end
            14'd7992 : begin out <= 64'b1010010100010110001010000010101100101010010000000010101000010100; end
            14'd7993 : begin out <= 64'b1010010101010101101010010100010010100001000011000010100111000110; end
            14'd7994 : begin out <= 64'b1010011001111010001010001011110010100011101101110010100100000100; end
            14'd7995 : begin out <= 64'b1010101110100110101001111010010100100001111011011010011010101110; end
            14'd7996 : begin out <= 64'b0010100010011000101000111100001110100110110001011010001101010001; end
            14'd7997 : begin out <= 64'b0010101010111110101010100101100010100110110011100001111110110110; end
            14'd7998 : begin out <= 64'b1010101101000000101010010000111100100111000010101010100111101010; end
            14'd7999 : begin out <= 64'b0010011111000111001000001010111010101010010000000010101101001111; end
            14'd8000 : begin out <= 64'b1010100001000000001010101110110010101011001110111010101101000110; end
            14'd8001 : begin out <= 64'b0010100010011101001010011011011100011000011001001010100100010100; end
            14'd8002 : begin out <= 64'b1010100100100000101010110001110010101010100111101010101100101100; end
            14'd8003 : begin out <= 64'b0010011101100011101010110010010110011001101001101010000001101000; end
            14'd8004 : begin out <= 64'b1010101101000100101010110000011000011000000001001010100000000011; end
            14'd8005 : begin out <= 64'b0001111011100111101001001111011100101001110001100001110100000010; end
            14'd8006 : begin out <= 64'b1001000101010111001010001001110000101010100010000010100010101001; end
            14'd8007 : begin out <= 64'b1010011001111000001001110110001010101011111010010010101000110100; end
            14'd8008 : begin out <= 64'b0010100101110010101010010000000100101000110001111010100000110010; end
            14'd8009 : begin out <= 64'b1001111101110000001010110101000110100010101100010010011101111100; end
            14'd8010 : begin out <= 64'b1001111100011110001010100110111110100111100000010010100000010110; end
            14'd8011 : begin out <= 64'b0010100101010000101000110100110000101000101010110010101111000001; end
            14'd8012 : begin out <= 64'b0010001100000001101000011100111100101001010111111010101100111111; end
            14'd8013 : begin out <= 64'b1010010100001100001010011010010010101000101110010010101101101000; end
            14'd8014 : begin out <= 64'b1001010000011000001010110111010010101010101110000010100111100100; end
            14'd8015 : begin out <= 64'b0010100111010000101000000001010000101010000001010010101001000101; end
            14'd8016 : begin out <= 64'b1010100010011100001001010110000100100001011110110010100011001001; end
            14'd8017 : begin out <= 64'b0010100100000101101010100101000110101001111110001010001101000101; end
            14'd8018 : begin out <= 64'b1001111111000011001010100010010100101011110001010010100110011000; end
            14'd8019 : begin out <= 64'b0010010101100101001010000100101010101001111000001010101000001100; end
            14'd8020 : begin out <= 64'b1001100000011001001010111100001000010100110001111010100010000010; end
            14'd8021 : begin out <= 64'b1010101101111110001010101111010100100100010010001010100000010100; end
            14'd8022 : begin out <= 64'b1010011010011001101010111011101110101000001101111010101010010001; end
            14'd8023 : begin out <= 64'b0010010000000001001010000011110110100110011001110010101110100100; end
            14'd8024 : begin out <= 64'b0010011111000010001010000100111110100110101111010010010000010000; end
            14'd8025 : begin out <= 64'b0010101001111011001001110110100100100101001110101010100110110100; end
            14'd8026 : begin out <= 64'b1010100110001000100100101001101100101010000010010010010101101111; end
            14'd8027 : begin out <= 64'b0001110110100010101010001000001110101011111001110010011111101000; end
            14'd8028 : begin out <= 64'b1010101100110101101010010000110000011010010001101010101100010001; end
            14'd8029 : begin out <= 64'b0010001001101000001010101010101110101011100100110010001001001100; end
            14'd8030 : begin out <= 64'b0010011010101110101010111101000100100101011111011010011000110100; end
            14'd8031 : begin out <= 64'b0010100101000010001010010010011000101010011000110001111000011101; end
            14'd8032 : begin out <= 64'b0010011011100110101001001001111110100101000000000010001100001000; end
            14'd8033 : begin out <= 64'b1010101101001010001001010001001000101011001010011001101011110011; end
            14'd8034 : begin out <= 64'b0010101110111000101010111110001100101000000110111010100101100110; end
            14'd8035 : begin out <= 64'b1001110100111011001010011010111010100100110101101010100010100001; end
            14'd8036 : begin out <= 64'b0010011001000000101010001011110000001110001101001010101101110111; end
            14'd8037 : begin out <= 64'b0010011110110000001010001011100000100000010100100010010001100101; end
            14'd8038 : begin out <= 64'b0010100101100001101001101001110000101011001010010001010100100100; end
            14'd8039 : begin out <= 64'b1010100111011111001000101001100010100001110001110010101011011111; end
            14'd8040 : begin out <= 64'b1010011111111001001001111010000000100110000010111010000011110100; end
            14'd8041 : begin out <= 64'b1010000110110101100110111001111100101001100010111010011100000010; end
            14'd8042 : begin out <= 64'b1001110011001101100111100001011100100010010011111010100000101000; end
            14'd8043 : begin out <= 64'b0010101011111010001010110110000010101000001001111010101010111100; end
            14'd8044 : begin out <= 64'b0010101111111100101001000000001000101011011010110001100010010000; end
            14'd8045 : begin out <= 64'b1010011100010111001010111011001110101001011000000010101011101101; end
            14'd8046 : begin out <= 64'b1010000111110010100111110111011010101001001100011010010100110010; end
            14'd8047 : begin out <= 64'b0010100011110100101000000111010010101001111000001010011111100100; end
            14'd8048 : begin out <= 64'b1010101110011100101001110010111100101011101010110010101001000011; end
            14'd8049 : begin out <= 64'b1010100100100011001000101000011110100101000000000010100001100011; end
            14'd8050 : begin out <= 64'b1010101011001010101010010010011000100110100000111010100000010110; end
            14'd8051 : begin out <= 64'b0010100111001010001010110100010010101001001010010010000000100100; end
            14'd8052 : begin out <= 64'b0010100110011000100111101011110100101011111101000010101110001110; end
            14'd8053 : begin out <= 64'b1010110000001000001001100010010000101100000010010010010010101111; end
            14'd8054 : begin out <= 64'b0010001111010100001001100011110010100010000011101010011111011111; end
            14'd8055 : begin out <= 64'b1010000101110100001010010011001010100101001110101010100010000101; end
            14'd8056 : begin out <= 64'b0010011110110111001010001110101010101010111001100010010010110101; end
            14'd8057 : begin out <= 64'b0010101111000001000110111101110000100100010100010010001110110100; end
            14'd8058 : begin out <= 64'b0010101000001000100110000000010000101000110001011001111011001010; end
            14'd8059 : begin out <= 64'b1010010011100000101001000011010010101000001001000010001111011110; end
            14'd8060 : begin out <= 64'b1010100011001101101001011011000000101001010110101010011010011100; end
            14'd8061 : begin out <= 64'b1010101111001001101000001010101110100010100101000010100010101100; end
            14'd8062 : begin out <= 64'b0010010011001101101010101110001000100101011010110010000000101011; end
            14'd8063 : begin out <= 64'b0010100111010100000111011111110110100101100110111010100101000010; end
            14'd8064 : begin out <= 64'b0010101101101011001010010110101010101000111011110010101111011001; end
            14'd8065 : begin out <= 64'b0010001110101111101010011000110010011110001010110001111000000000; end
            14'd8066 : begin out <= 64'b1010101000011011000010100110111000101010000001110001111001100000; end
            14'd8067 : begin out <= 64'b0000111011100000001001101101111100100101000101000010110000000110; end
            14'd8068 : begin out <= 64'b0010010101010000101010001100110110100100010111011010010101000010; end
            14'd8069 : begin out <= 64'b1010100010000101101001100001100010101001101001010010010000001100; end
            14'd8070 : begin out <= 64'b0010011000100101101010011010111010101011100001110010101000010010; end
            14'd8071 : begin out <= 64'b1010100101000011100111110001010010100110010101011010100010010010; end
            14'd8072 : begin out <= 64'b0010100111101101001001101111000100100111101011101010100010100000; end
            14'd8073 : begin out <= 64'b1010001001001010101000111010111100100110111100100001101101001010; end
            14'd8074 : begin out <= 64'b0001100010110011101000001011110000100011100100110010100010110100; end
            14'd8075 : begin out <= 64'b0010100101011111101001011111101110101011010100100001110111001001; end
            14'd8076 : begin out <= 64'b1010100010010110101010011110111100100000011110001010011110100101; end
            14'd8077 : begin out <= 64'b1010000000110111001010101011101010101001011010101010010010000000; end
            14'd8078 : begin out <= 64'b1010100110010101101001111001000000101001010101010010100100010000; end
            14'd8079 : begin out <= 64'b1010010110010110101000011001100000101001110000001010100110001100; end
            14'd8080 : begin out <= 64'b0001110111101010001001100001001100101001100001101010011010101000; end
            14'd8081 : begin out <= 64'b0010000111011000101010000000101110011110110111100010000100101101; end
            14'd8082 : begin out <= 64'b1010010011100101101010101101001010101011110100111010101110010111; end
            14'd8083 : begin out <= 64'b0010000011000110101010101000110110101010101110010010100010011110; end
            14'd8084 : begin out <= 64'b0010100001010011101001011000101110101011001100110010101101100000; end
            14'd8085 : begin out <= 64'b1010101011010000101001001111011000101010101110101010101001101110; end
            14'd8086 : begin out <= 64'b1010100000001100001010111101100100101010000111101010010110111001; end
            14'd8087 : begin out <= 64'b1010001110010001101001110010100010101000101100011010100100101000; end
            14'd8088 : begin out <= 64'b0010011111000110000110001101101000101001101001001010001111000101; end
            14'd8089 : begin out <= 64'b1010101111100110101001001101001100101001100100011010100010101111; end
            14'd8090 : begin out <= 64'b1010011011011100001010110100010010101010101101001010100010010010; end
            14'd8091 : begin out <= 64'b0010000001110110001010010101111100100001110000001010010100000111; end
            14'd8092 : begin out <= 64'b1010101000111001001010110110101010101001000000000010100110100100; end
            14'd8093 : begin out <= 64'b1010101110111000000111001100100110011111001001010010101001011001; end
            14'd8094 : begin out <= 64'b0001111011001110101000001101101000100001011111000010110001001010; end
            14'd8095 : begin out <= 64'b1010011101100010001001010001011100100101001101110010100010010101; end
            14'd8096 : begin out <= 64'b1010011011100110101010001101001010100011100111111010101010000101; end
            14'd8097 : begin out <= 64'b0001110010001101001010010011011100100101101101111001101000101110; end
            14'd8098 : begin out <= 64'b1010101000101000101010100111111100101011001010111010100010001100; end
            14'd8099 : begin out <= 64'b1010010001001100101000111010001010010101100100001010101011111110; end
            14'd8100 : begin out <= 64'b0010100001110111101001010000011010011111101001001010100100000111; end
            14'd8101 : begin out <= 64'b1010101011001001100111111110000010100000110000000010001010110000; end
            14'd8102 : begin out <= 64'b1010011000011100000111110001001000100111111111101010010100010101; end
            14'd8103 : begin out <= 64'b0010100110001001101000110100011010101010000101111010110000110111; end
            14'd8104 : begin out <= 64'b0010000101010110001000110011111110100001111101101010011010011111; end
            14'd8105 : begin out <= 64'b0001100110001110101001001000001100101001111101110010100011010000; end
            14'd8106 : begin out <= 64'b0010101010110101001010001010111100101000111011001010010001001110; end
            14'd8107 : begin out <= 64'b0010001010111001000010100011001010101011111001010010101101011010; end
            14'd8108 : begin out <= 64'b1001111100000110001001110010000000101011100000000010010010010010; end
            14'd8109 : begin out <= 64'b1010101110010011101010010111100000100111111101110010101100110110; end
            14'd8110 : begin out <= 64'b0001101011010011001010010000101100101000110100100010010100101011; end
            14'd8111 : begin out <= 64'b0010011100100111101000001010111000100101110101111010100011000011; end
            14'd8112 : begin out <= 64'b0010101011100000001000101100010000101000111011100010101001101011; end
            14'd8113 : begin out <= 64'b0010101010011110100111010101010000101010001000100010101011101011; end
            14'd8114 : begin out <= 64'b1010011001010100101010111110001000100001000010100010100111001011; end
            14'd8115 : begin out <= 64'b0010010011011100101000101100001010011101001110000010100001101010; end
            14'd8116 : begin out <= 64'b0010101101000000001010101101001100101010110110010010101000101010; end
            14'd8117 : begin out <= 64'b0010001001110010101001111000101100100110101100001010100010001000; end
            14'd8118 : begin out <= 64'b0010100000000001101010101010110010100110011000101001111110100001; end
            14'd8119 : begin out <= 64'b0010100001011100101001011011010110101010001010001010011011101000; end
            14'd8120 : begin out <= 64'b1001111111001001101010100100010010101100001100011010001110011011; end
            14'd8121 : begin out <= 64'b1010101011100100101010001111111000101011110000100010101010110001; end
            14'd8122 : begin out <= 64'b1010100011111010001010011110010110010110000111110010011100100001; end
            14'd8123 : begin out <= 64'b0001110100100101001001011100000100100110100000000010100010011100; end
            14'd8124 : begin out <= 64'b1010000100001011101000000100101000011100111110010010000011110101; end
            14'd8125 : begin out <= 64'b0010010100101110101010011010100110101001111010001010000111001101; end
            14'd8126 : begin out <= 64'b0010001101100011101010010100011000100110010001110010101010111101; end
            14'd8127 : begin out <= 64'b0010101001101100100111100010001100011011001111110010100001001000; end
            14'd8128 : begin out <= 64'b0001111011000001001010011111111100101000110001011010011011111011; end
            14'd8129 : begin out <= 64'b0010100010110000001010111011000000100110100000110001101110000100; end
            14'd8130 : begin out <= 64'b1010100110001011001010000110001010100101100001101010100111101110; end
            14'd8131 : begin out <= 64'b0010000111000110001010000101001100100001101001000010100110110110; end
            14'd8132 : begin out <= 64'b1010010011111110101001010000110110011000100010001010100100001111; end
            14'd8133 : begin out <= 64'b1010010000011010101010011010110110011100101110100010000001011110; end
            14'd8134 : begin out <= 64'b0010010101110100001001101010000000101000001100110010101000011000; end
            14'd8135 : begin out <= 64'b0010101000100100001010101101110100100111100001001010000110011010; end
            14'd8136 : begin out <= 64'b0010101000100110001010001100100010101000100111010010101011111000; end
            14'd8137 : begin out <= 64'b0010100110100001001000001111100000101010110101101010010111001110; end
            14'd8138 : begin out <= 64'b1010101110110101001010000011001010100000010101110010100110111010; end
            14'd8139 : begin out <= 64'b1010100100000110001000101001010100100101101111011010000010011010; end
            14'd8140 : begin out <= 64'b0010000001011010100000111101011000011001011000001010100100100100; end
            14'd8141 : begin out <= 64'b1010011010000111001010100010111010100100001011000010000111000000; end
            14'd8142 : begin out <= 64'b0010000010010110001010101101001000101011010111001010000101001011; end
            14'd8143 : begin out <= 64'b1010010001011000101001011111101100100000000101011010011000010010; end
            14'd8144 : begin out <= 64'b0010100110010000100101111100101010011011000001000010101100011001; end
            14'd8145 : begin out <= 64'b0010001101010110101010110100011100101011011010100010011100010011; end
            14'd8146 : begin out <= 64'b1010011100100101000111111110010110100100011110000000101101110111; end
            14'd8147 : begin out <= 64'b1010010101100010101001000010001100011110111010111010110000010011; end
            14'd8148 : begin out <= 64'b1010101010110100001010010100111100101011111000010010010010101110; end
            14'd8149 : begin out <= 64'b1010011001110010100100110110100100100000001001111010100111111000; end
            14'd8150 : begin out <= 64'b1010101110011110100111011101010000101000010101111010011000000101; end
            14'd8151 : begin out <= 64'b0010100101101100101010111100110000101001100001001010100111010111; end
            14'd8152 : begin out <= 64'b1010101001011100100111110010001010101011001100100010101100010001; end
            14'd8153 : begin out <= 64'b1010011010001100101001011010010100101000101011101010011011101001; end
            14'd8154 : begin out <= 64'b1010101101110101101001010100001010101011101110000010001111010011; end
            14'd8155 : begin out <= 64'b1010101000101011001001010010010010101011000011010010100011111101; end
            14'd8156 : begin out <= 64'b0010011101111011101001001010001100101000101001011010101100100001; end
            14'd8157 : begin out <= 64'b0010011001011001101010110110011010100001010010100010101100000100; end
            14'd8158 : begin out <= 64'b1010000110110001101010000010100010101011101010000010011010001110; end
            14'd8159 : begin out <= 64'b0001111000011101100001010000010000100111011100001010001011111001; end
            14'd8160 : begin out <= 64'b1010100101010001101010001000100000100101000001001000000000011111; end
            14'd8161 : begin out <= 64'b0010101100011110101010111010010010100110000100101010100011000101; end
            14'd8162 : begin out <= 64'b0010110000000100101001111110110000011011110001101010001010010010; end
            14'd8163 : begin out <= 64'b1010101011000110101010000111010110101001110111011001110101101010; end
            14'd8164 : begin out <= 64'b0010010101010011001010100111001010010000111011011010100110011000; end
            14'd8165 : begin out <= 64'b1010100001010001100011111010011000101000011001000001100111000111; end
            14'd8166 : begin out <= 64'b1001111110101011001001010111110000101000011001110010000001101000; end
            14'd8167 : begin out <= 64'b1001111011110100101010100010110100100111101101111010001010111000; end
            14'd8168 : begin out <= 64'b0010100001001011101010001100000000100100000100110010101010100110; end
            14'd8169 : begin out <= 64'b1010101100111100101010101000011010100010011011001010010011010010; end
            14'd8170 : begin out <= 64'b1010010111001000001010000110101100100100001000010001001000110101; end
            14'd8171 : begin out <= 64'b0001111010110010101001100010111010101000011011100010000100011110; end
            14'd8172 : begin out <= 64'b1010101001111111101010100010100100100110100011011010000111000101; end
            14'd8173 : begin out <= 64'b1010010100001100001010100011010000101010101000000010010001110001; end
            14'd8174 : begin out <= 64'b1010100001011100001000100101000110011111110111010001111111000111; end
            14'd8175 : begin out <= 64'b1010100000011110101010000111011100101000001111011001111110000100; end
            14'd8176 : begin out <= 64'b0010100011100000001001111010011110011101110001000010100111000000; end
            14'd8177 : begin out <= 64'b1001100101110100101010101001000010101010110101111010010010101110; end
            14'd8178 : begin out <= 64'b0010011110101100101001110110000100100011100110110010100001001000; end
            14'd8179 : begin out <= 64'b0010001110011111101001110001000000100100000101000010101001101111; end
            14'd8180 : begin out <= 64'b0010011111111000101010010100100010101000000100111010100101100101; end
            14'd8181 : begin out <= 64'b1010100110001010001010101111101010101000001010101010010101101000; end
            14'd8182 : begin out <= 64'b1010101010010011101010000001010110101001000111000010011110011101; end
            14'd8183 : begin out <= 64'b1010010110011101101010100000010100101001100000111010101001000000; end
            14'd8184 : begin out <= 64'b1010101101011110001010000011010000100010000111001010101000100000; end
            14'd8185 : begin out <= 64'b0010101110001001101010111000101000100110110010100010110000101110; end
            14'd8186 : begin out <= 64'b1010001100101111101010111011100000011011100000101010110001110010; end
            14'd8187 : begin out <= 64'b0010100111000001001001000010111010100010001010010010010110011010; end
            14'd8188 : begin out <= 64'b1010010100111101101001001001100000011101101110010010010011100111; end
            14'd8189 : begin out <= 64'b0010101011000011001000100101101000011100111011101010100110010001; end
            14'd8190 : begin out <= 64'b1010011001100111001010111100101010101010010000110010100101000011; end
            14'd8191 : begin out <= 64'b1010100100110010001001001101000000011000011000110010100000000100; end
            14'd8192 : begin out <= 64'b1010101000011100101000000011110110101001110001111010100100100110; end
            14'd8193 : begin out <= 64'b0010100111001100101011000000001100100111100110001010100110111111; end
            14'd8194 : begin out <= 64'b1010011010010010101001111111110010100100001111111010010111001101; end
            14'd8195 : begin out <= 64'b0010000101111111001000010110010010101000100011111010000001011110; end
            14'd8196 : begin out <= 64'b1010100010000000100111111001110100101001000001110010101101001001; end
            14'd8197 : begin out <= 64'b1010000111011101100111110111111000001101100000001010100101111001; end
            14'd8198 : begin out <= 64'b0001110110100100000111111011001100101010000110110010011110111110; end
            14'd8199 : begin out <= 64'b0010101000111000101010101001110100101011100100110010100101100110; end
            14'd8200 : begin out <= 64'b0010101011100001100111101001010000100011010000101010101100110000; end
            14'd8201 : begin out <= 64'b0010100011101111001010010101110100101011001101111010010010111101; end
            14'd8202 : begin out <= 64'b0001110001101000000111000110011010101001100100101010101101110000; end
            14'd8203 : begin out <= 64'b0010010101000000001010110010011000101001001010001001111000011000; end
            14'd8204 : begin out <= 64'b0010001001011010001001110110000100101011101000110001110110111000; end
            14'd8205 : begin out <= 64'b0010100000101110101010001101010000010001000111111010100101010001; end
            14'd8206 : begin out <= 64'b0010011101111110001001000100000100101001100010010010101000001110; end
            14'd8207 : begin out <= 64'b1010100110111110001010101101001000101001110110110010000000101001; end
            14'd8208 : begin out <= 64'b0010101111101000101001101111011010101010001010101010010111010111; end
            14'd8209 : begin out <= 64'b1010101110010001101011000101000010101001110001011010101010111001; end
            14'd8210 : begin out <= 64'b0010010010101111101001111011001000101000000110001010010101000110; end
            14'd8211 : begin out <= 64'b0010101110010001101001000110000000101000100010000010000001001000; end
            14'd8212 : begin out <= 64'b0010100010100000001000110110111010101000100110011010101100100111; end
            14'd8213 : begin out <= 64'b0010100010100101101010000111010010100000011000101010101111110001; end
            14'd8214 : begin out <= 64'b0010100101111010001001010110101110100110010010100010011101001110; end
            14'd8215 : begin out <= 64'b1010100011010100101001010010101010101000011100101010101110011110; end
            14'd8216 : begin out <= 64'b0010010111010110101010001101011100100100001110101010101001100110; end
            14'd8217 : begin out <= 64'b1010010111100111001000010011000110100110100001010010101100011100; end
            14'd8218 : begin out <= 64'b0010010011000001001001111011010100101010111010001001110110101011; end
            14'd8219 : begin out <= 64'b1010010001101111101010010100001000100111001000010010010001001000; end
            14'd8220 : begin out <= 64'b0010010101110110000111001110001010101011111101110010011110011010; end
            14'd8221 : begin out <= 64'b1010000010100001000110100101100100101000100001111010100010100100; end
            14'd8222 : begin out <= 64'b0001110101001100101001001111011100100111001001100001000100000010; end
            14'd8223 : begin out <= 64'b0010011000011110101010101101000010100100001010100010100011001010; end
            14'd8224 : begin out <= 64'b0010000110010101100011000101111010101000101011101010100011010010; end
            14'd8225 : begin out <= 64'b0010101110010110101001101001100010101010001011001001100001101010; end
            14'd8226 : begin out <= 64'b1010011101000111101010110000111010100100111111000010010011001100; end
            14'd8227 : begin out <= 64'b0010100010100110101010011100101100100111010001101010010010001110; end
            14'd8228 : begin out <= 64'b1010011101101100001000101111010100100110011101101010011101111010; end
            14'd8229 : begin out <= 64'b0010000100010000101010110111101010100000110001010001110011101001; end
            14'd8230 : begin out <= 64'b1010100111100111101000000010101000100110010010000010000010010101; end
            14'd8231 : begin out <= 64'b1010101010000001101000001111110010101000101000110010010101010010; end
            14'd8232 : begin out <= 64'b0010001110101011001001101110100000100011100010110010010001110000; end
            14'd8233 : begin out <= 64'b1001111010001110001000011101001010100111010001011010100111010010; end
            14'd8234 : begin out <= 64'b0010101001100011001001010001000100100101000111111010100000010111; end
            14'd8235 : begin out <= 64'b0001110101001010001001010001110110100100001010110001001100101111; end
            14'd8236 : begin out <= 64'b1010100010000101101000011010010110100010101010011010101010001111; end
            14'd8237 : begin out <= 64'b1010101000101110101010000100001100100111001101110010001111010011; end
            14'd8238 : begin out <= 64'b1010010110011110000100011001000000101010001011111010101101011001; end
            14'd8239 : begin out <= 64'b1010011011100001101001001011110010100101010000001010000110011010; end
            14'd8240 : begin out <= 64'b1010101100101000101010111101100000101011000011110010011000010010; end
            14'd8241 : begin out <= 64'b0010101000010111001010100010001110101000010111010010010001011100; end
            14'd8242 : begin out <= 64'b0010100101001010001010000111111010100110100010000010100011110000; end
            14'd8243 : begin out <= 64'b1010101110010101101000000101110100101011011110000010101110010011; end
            14'd8244 : begin out <= 64'b1010011000110011000111001110101110100100010001011010001111000000; end
            14'd8245 : begin out <= 64'b0010101010100110001000011100101000101010001100000010010000011001; end
            14'd8246 : begin out <= 64'b1001111101101101000110100111101100100100001001101010010100101111; end
            14'd8247 : begin out <= 64'b0010010000010110001010000010101010101001010100110010101010001111; end
            14'd8248 : begin out <= 64'b1001110111000010000110111011011100100010001100001010100101011011; end
            14'd8249 : begin out <= 64'b1010100001001101101001011001001000100111001111101010100111101110; end
            14'd8250 : begin out <= 64'b0010100100000111101000111001010010100000101101011010000101110110; end
            14'd8251 : begin out <= 64'b0001011101110001100101010011110110101010111111000010001011100000; end
            14'd8252 : begin out <= 64'b1010101000101010001001011001101000100011010000111010010101010100; end
            14'd8253 : begin out <= 64'b1010101001101101101001110000101110101011111001011010100010001011; end
            14'd8254 : begin out <= 64'b0010101100111111000111011100001010011100001111100010011000110011; end
            14'd8255 : begin out <= 64'b1010101101001110101010110110011110100110001110101010101011100110; end
            14'd8256 : begin out <= 64'b0010101110000110100110001110010000100011111100100010101100101011; end
            14'd8257 : begin out <= 64'b1010100110101010001010101111101110101001001110011010001010010101; end
            14'd8258 : begin out <= 64'b1010101001100110101010001100111000101010011000100010101100111100; end
            14'd8259 : begin out <= 64'b1010100111111111001000000101010010101011001110001010101000010000; end
            14'd8260 : begin out <= 64'b1001101111100000001001101110100110011100110011010010101001010001; end
            14'd8261 : begin out <= 64'b1010101101110111101010101011001110100110000100111010101100110010; end
            14'd8262 : begin out <= 64'b1010010110011011001000110111011100100101111101101010010100011010; end
            14'd8263 : begin out <= 64'b1010011011100011101010010100011100100010001111011001011110101100; end
            14'd8264 : begin out <= 64'b0001110110100001001010000101001000011101101011110010001100000010; end
            14'd8265 : begin out <= 64'b0010010000110101101000000011100010100011000100110010101111000010; end
            14'd8266 : begin out <= 64'b1010101101101101101011000010111110101000011111000010010011001011; end
            14'd8267 : begin out <= 64'b0010100100111100101010101001110000100111100111001010100111001101; end
            14'd8268 : begin out <= 64'b1010011011010101101001011010001010100001001001110010100110110111; end
            14'd8269 : begin out <= 64'b0001011010011000101010110001110000101011001100010001100110100110; end
            14'd8270 : begin out <= 64'b0010100101100010101000100111101000100101011101000001111010111101; end
            14'd8271 : begin out <= 64'b0001111100000110101010011100100000101011110111100001100100111010; end
            14'd8272 : begin out <= 64'b0010100111001110101001001110101000101000010011111001110010100101; end
            14'd8273 : begin out <= 64'b0010100111100111000110010100111100010101010000100010000001011110; end
            14'd8274 : begin out <= 64'b1000100100110010100101010011101110101000010000001000111010101111; end
            14'd8275 : begin out <= 64'b1010101100110000101011000101010100100100110110111010101110100101; end
            14'd8276 : begin out <= 64'b1001110011000001001001111011001100101001011010000010100001110101; end
            14'd8277 : begin out <= 64'b1010100010011101101001111001101110101000101111111010010110001100; end
            14'd8278 : begin out <= 64'b1010101111000101001000100011100100100010111101110010101010111010; end
            14'd8279 : begin out <= 64'b0010100111100101001010001000010100101010011101111010101100011010; end
            14'd8280 : begin out <= 64'b1010011101110001001001001011010100100101100000010010100111111010; end
            14'd8281 : begin out <= 64'b1010110000001000001000000000100010100110010101101010010011010010; end
            14'd8282 : begin out <= 64'b1001100101111000101010100101111010011100100111000010100101000111; end
            14'd8283 : begin out <= 64'b1001111100111011001010110100000000101011100000001001110101011111; end
            14'd8284 : begin out <= 64'b0001110010110110001010010010111000100111111101011010000011001111; end
            14'd8285 : begin out <= 64'b1001011011100111001010110000101100101001111011010010101011001001; end
            14'd8286 : begin out <= 64'b0010100110010110001000111011101010101011011101111010100000110011; end
            14'd8287 : begin out <= 64'b0001110110000010001010011101001000101000111011011001010011011100; end
            14'd8288 : begin out <= 64'b0010011001100010100100110100011010101001011010010010101000110101; end
            14'd8289 : begin out <= 64'b0010100110011101101001101110001110100100011011101010010010101001; end
            14'd8290 : begin out <= 64'b1010100011110011001001010010111100101011110111100010101010111111; end
            14'd8291 : begin out <= 64'b1010101110110101001000011110010000100111011010001010101010101011; end
            14'd8292 : begin out <= 64'b0010100011111010001001110010101100100000011110110010011001101010; end
            14'd8293 : begin out <= 64'b0010101010111100101010110100111110100110001111010010010110100101; end
            14'd8294 : begin out <= 64'b1010101011110001001000000111010000101000100010110010101101111011; end
            14'd8295 : begin out <= 64'b0010010010110101000111011111111000100011111000000001100110100101; end
            14'd8296 : begin out <= 64'b0010101100001100101001001011001010101011110010110010101111011111; end
            14'd8297 : begin out <= 64'b1010010001111101101010110001100110101011001001011010100001001010; end
            14'd8298 : begin out <= 64'b0010100001001001101000111110101100100101111110001010100001100000; end
            14'd8299 : begin out <= 64'b1010010001011111001000111011000010100100011110110010100000110100; end
            14'd8300 : begin out <= 64'b0010100110100001101000010110110010101010011011110010101111100101; end
            14'd8301 : begin out <= 64'b1010000001001000101010010001111010100101110000100010011101101100; end
            14'd8302 : begin out <= 64'b1010010010011001001010111101000000101010001110010010011010010001; end
            14'd8303 : begin out <= 64'b1010011101100010001010000000101100101010001000000001110001001011; end
            14'd8304 : begin out <= 64'b1001010100100101101010011011000110101010011100100010100001011101; end
            14'd8305 : begin out <= 64'b1001110011110101101000000011101110100100111101011010100100101100; end
            14'd8306 : begin out <= 64'b0010101011010010001000011110001110101011110111010010011000000010; end
            14'd8307 : begin out <= 64'b1010000100000011101000001110110010011110010011010010100001011010; end
            14'd8308 : begin out <= 64'b1010100100011000001010111010101010101001100100111010100111010100; end
            14'd8309 : begin out <= 64'b0010101101000101101010000110010010100110101100101010100110001001; end
            14'd8310 : begin out <= 64'b1010101000101110101000100110001110100011111100001010010010111101; end
            14'd8311 : begin out <= 64'b1010101000101010101010101011101000100100101010001001011001111001; end
            14'd8312 : begin out <= 64'b1010010011101101101001111100111100101011000110110010101010100110; end
            14'd8313 : begin out <= 64'b0010100001011001001010001111100100011101000111110010011000101110; end
            14'd8314 : begin out <= 64'b0010011101101000101000110011000000101011001001000010101010011000; end
            14'd8315 : begin out <= 64'b0010010100110001001010111010000110101001010001010001101110001110; end
            14'd8316 : begin out <= 64'b0010100000001100101010011000010010011100100111110010100000010010; end
            14'd8317 : begin out <= 64'b1010100111000110001000001111101110101010001110011010100010111000; end
            14'd8318 : begin out <= 64'b0010101110010000101001100000000000101000111101100010000110011100; end
            14'd8319 : begin out <= 64'b1010100011010110101011000100100100100110111000100010011010101010; end
            14'd8320 : begin out <= 64'b1010010100011110101010101011100010011111100000100010010000100011; end
            14'd8321 : begin out <= 64'b0010100010001000000110011111001010100101101010010010100011000011; end
            14'd8322 : begin out <= 64'b0010101100010010001010001100101000101010000001110010100101011111; end
            14'd8323 : begin out <= 64'b1010100111001001101000010001110110101011110100010010101011100011; end
            14'd8324 : begin out <= 64'b1000110101101010101010100110101010101011001101101010001011111001; end
            14'd8325 : begin out <= 64'b1010010010000010101010011101011100100111111010110010100001001100; end
            14'd8326 : begin out <= 64'b0010011000011101001011000110101100101010011100000010101101101100; end
            14'd8327 : begin out <= 64'b0010101111110001101000011000100010100111011001001010101100001110; end
            14'd8328 : begin out <= 64'b0010011111101011001010100001101000100111101000011010100010110000; end
            14'd8329 : begin out <= 64'b1010100001011101001000100010001010101000111000011010001100001101; end
            14'd8330 : begin out <= 64'b1010011001111111101000001001000100011110100000110001100111101010; end
            14'd8331 : begin out <= 64'b1001101000000111101010011110111110101000000001100010100010101011; end
            14'd8332 : begin out <= 64'b1010011111011101101001011001101100101001011100011010100101010101; end
            14'd8333 : begin out <= 64'b0010011111111101101001000000001000101000111001100010100101010010; end
            14'd8334 : begin out <= 64'b0010101101101010101001110011001000100101101101101010100111011000; end
            14'd8335 : begin out <= 64'b1001111100010000101010110111010110101011100010101010010110100011; end
            14'd8336 : begin out <= 64'b0010101001010100100111010010000010101000101100101010100010010100; end
            14'd8337 : begin out <= 64'b0010000001011010001010000011001000101011001010110010100101000000; end
            14'd8338 : begin out <= 64'b1010101001100101101000100001001100101010010101000010100111111000; end
            14'd8339 : begin out <= 64'b0010101111000011101001101110111010100010011110110010101000011001; end
            14'd8340 : begin out <= 64'b1010011011010001001000001111100110101000001110101010101110110001; end
            14'd8341 : begin out <= 64'b0010101111101011101000000011111110100110101101111010100110010110; end
            14'd8342 : begin out <= 64'b0001111110111110101001011110011010011100010000111010101101111101; end
            14'd8343 : begin out <= 64'b1010101100011111001001000110000100100110000110010010011010100110; end
            14'd8344 : begin out <= 64'b1010100010010011101010100011000000101001111011100010010101100101; end
            14'd8345 : begin out <= 64'b0010101101000100001001101111010010100111001100011010011111111111; end
            14'd8346 : begin out <= 64'b0010101011101101101010011101000110100101111011100010101110110110; end
            14'd8347 : begin out <= 64'b0010101110101011001010001001000000101011011101010010011011110110; end
            14'd8348 : begin out <= 64'b1010010111111100000100111110011010011101101000110010100001111101; end
            14'd8349 : begin out <= 64'b0010010001010001001000010010000110100101111000011010101111000101; end
            14'd8350 : begin out <= 64'b1001011100001000101001100110010000101000101101011010010110000100; end
            14'd8351 : begin out <= 64'b1010000001001101001000101110110100101010011110010010010110101101; end
            14'd8352 : begin out <= 64'b1001110011011111101010010000100000101010100100011010101100000000; end
            14'd8353 : begin out <= 64'b0000000011110100101010101011010010101011011101010010101110001010; end
            14'd8354 : begin out <= 64'b1010100100110011001010000110010010100100110001100010010101101011; end
            14'd8355 : begin out <= 64'b0010000100010000001010001100111000101011011000111010011001001111; end
            14'd8356 : begin out <= 64'b1010011001001110101010011011111100101010001100010010100000101010; end
            14'd8357 : begin out <= 64'b1010101001001011101010001001110110100111011101100001110100100010; end
            14'd8358 : begin out <= 64'b1001100101001001101010011100000000100101100001110010101110100011; end
            14'd8359 : begin out <= 64'b0001100000010010001010000011101100011001000010101001111000111001; end
            14'd8360 : begin out <= 64'b1010010101001110101000100011100010101001110100100010100111111001; end
            14'd8361 : begin out <= 64'b1010001000010000100111100011000000101010001101000010010111101001; end
            14'd8362 : begin out <= 64'b0010101100001111101000111100101110101011100110101010000100111000; end
            14'd8363 : begin out <= 64'b1010011010001010001010010100011010101010111001101010100100000001; end
            14'd8364 : begin out <= 64'b0010101011110100101000101011001000101010010111101010101111010111; end
            14'd8365 : begin out <= 64'b1010100110110000101001011011110100100000111111000010101010100111; end
            14'd8366 : begin out <= 64'b1001101000100011000111111010010000101001000111110010100000111101; end
            14'd8367 : begin out <= 64'b0010101001110101001001000101010010101010110000101010000001010000; end
            14'd8368 : begin out <= 64'b0010011101010101101010000011101100100001001110001010101100110100; end
            14'd8369 : begin out <= 64'b0001100110110111000101111010011010101001001101000010010011111110; end
            14'd8370 : begin out <= 64'b0010001010110010001010101110100000100001100101000010100110100100; end
            14'd8371 : begin out <= 64'b0010010010100111001001001100011000101100000000000010100111101001; end
            14'd8372 : begin out <= 64'b1001010110000101001000111010101000101010000010100010000001101010; end
            14'd8373 : begin out <= 64'b0010010011100110001010001111001100101000011011100010011101010001; end
            14'd8374 : begin out <= 64'b0010011011100000001001110110110000101010010101010010101010000010; end
            14'd8375 : begin out <= 64'b1010100100000100001010010000110110101001111101010010100001011011; end
            14'd8376 : begin out <= 64'b0001111110001110001010101010100100101000000101101010001100000011; end
            14'd8377 : begin out <= 64'b0010001101000111101001111111100100101001100111001010011100011001; end
            14'd8378 : begin out <= 64'b1010011111101111101001101001100010100100100110010010100001110010; end
            14'd8379 : begin out <= 64'b1010100101110011001011000111000100101000110111110001000010001010; end
            14'd8380 : begin out <= 64'b1010010010111001101010010011000000101011110000010010000010110000; end
            14'd8381 : begin out <= 64'b1001101110100010100111111001101100100111000101111010100101011010; end
            14'd8382 : begin out <= 64'b1010011100001100101001001100111000101011001110010001111100110001; end
            14'd8383 : begin out <= 64'b1010001001000001101010110000110010011100000110111010101110110010; end
            14'd8384 : begin out <= 64'b0010000101001101000110010000011110101011100010010010100010101100; end
            14'd8385 : begin out <= 64'b1010001011001111001010011110110000101011100010101010101110011001; end
            14'd8386 : begin out <= 64'b1001111101101100001001101111001000011101111010011010101110000010; end
            14'd8387 : begin out <= 64'b0010101011101110101010000010111000101010110101101010010100000101; end
            14'd8388 : begin out <= 64'b1010011111001111101010011010001100101010110000010010100101000001; end
            14'd8389 : begin out <= 64'b1010101000001011101010001010001100101000000010101001101110001101; end
            14'd8390 : begin out <= 64'b1010100111111001000111000011110010100110101000000010000010100001; end
            14'd8391 : begin out <= 64'b0010100010100101001001000100111010100101010011101010000001011010; end
            14'd8392 : begin out <= 64'b0010100011110010101001001011001110101011111110010010010000011101; end
            14'd8393 : begin out <= 64'b0010010100000110101001000001101010101001100001101010101000000000; end
            14'd8394 : begin out <= 64'b0010100010011100101000001111111010100011000101100010101011011001; end
            14'd8395 : begin out <= 64'b1001111101111011001010011011001010011000111101101001111001111110; end
            14'd8396 : begin out <= 64'b1010100011101000001001100001111110101001001111001001010100110100; end
            14'd8397 : begin out <= 64'b1001110111110011001010001101110110100111001100001010101110111010; end
            14'd8398 : begin out <= 64'b0000101000101011101010010011011000101011110000000010101010010111; end
            14'd8399 : begin out <= 64'b0010101001110010001001010110010100101000101011111010101101101001; end
            14'd8400 : begin out <= 64'b0010101100100111001010110010001110100111001110011001010001111100; end
            14'd8401 : begin out <= 64'b1010010101110001001010001010001110101000101001000010000011100000; end
            14'd8402 : begin out <= 64'b1001111010101111101010010101111000100100010111000010001001010101; end
            14'd8403 : begin out <= 64'b1010101011111111000110111000111110100111100100111010101001110000; end
            14'd8404 : begin out <= 64'b1010101000010101001010001100010110101010010100001001011111010011; end
            14'd8405 : begin out <= 64'b0010011000101100001010110100101110101000101011001001100010000110; end
            14'd8406 : begin out <= 64'b1010101010001110101001110100001010011001110111101010010111100010; end
            14'd8407 : begin out <= 64'b1010000101110111101010011111111010100001101100100010101111011011; end
            14'd8408 : begin out <= 64'b1010101010001100101001011001111010101001000001000010001111010010; end
            14'd8409 : begin out <= 64'b0010011101110001101010011110001000100101011101101010100011001000; end
            14'd8410 : begin out <= 64'b0010000101111001001010010100000100101010011010100010010001100000; end
            14'd8411 : begin out <= 64'b0010101010000010101001000001110100101001101010110010100101010011; end
            14'd8412 : begin out <= 64'b0010100001011000101000000110000010101010111100111010100100010100; end
            14'd8413 : begin out <= 64'b1001110110000011101010000010001010101010111011111010100011010010; end
            14'd8414 : begin out <= 64'b1010010100001011000110111101011010100101100000110010101011010101; end
            14'd8415 : begin out <= 64'b0010101001111100101000000101110110101011101001110010100110101110; end
            14'd8416 : begin out <= 64'b0010101010011000101010111000101100101000100011100010010101100011; end
            14'd8417 : begin out <= 64'b0001110011000110000100101001000100100000100100011010011010001101; end
            14'd8418 : begin out <= 64'b1010100000110001101010010011010100101000110110101010100110011100; end
            14'd8419 : begin out <= 64'b0010100110011101101010001111101100101000010011001010101101011110; end
            14'd8420 : begin out <= 64'b0010010010001011001001111111000000101011111100001010010010111110; end
            14'd8421 : begin out <= 64'b1010101000111100101001100000011000101010001111110010010000110011; end
            14'd8422 : begin out <= 64'b0001001011011101001010011010101100100110100100111010101011110111; end
            14'd8423 : begin out <= 64'b0010101110101101001010000011110000101001000110100010100100011011; end
            14'd8424 : begin out <= 64'b0001111011000111101010101100001000101010100011111001110110101011; end
            14'd8425 : begin out <= 64'b1010001000001110101010100010111100011100110000100001111011100000; end
            14'd8426 : begin out <= 64'b0010101011000111001010001010010110101000111000111001110011111101; end
            14'd8427 : begin out <= 64'b1010100010110001101010001101001100100101111001100010101000110000; end
            14'd8428 : begin out <= 64'b0001110000111000001010011111010110100110110001010010101000001010; end
            14'd8429 : begin out <= 64'b0010100100100010001001111000100110100011111101100010101001100100; end
            14'd8430 : begin out <= 64'b0010101101011101101001110111100100101001101011001010010011011111; end
            14'd8431 : begin out <= 64'b0010101001001000001010100010110000101000000001111010101011010110; end
            14'd8432 : begin out <= 64'b1010101101100010001010100101011110101011001001101010101000000110; end
            14'd8433 : begin out <= 64'b0010100100011101001010000111100100100111110010110010100001111100; end
            14'd8434 : begin out <= 64'b1010101100101111101010001011001110011110100001000010000111111010; end
            14'd8435 : begin out <= 64'b0010001010111110101000111111011100100110001000101010100000111001; end
            14'd8436 : begin out <= 64'b0010100010011101101010011010110010100000110000000010101101111110; end
            14'd8437 : begin out <= 64'b1000100001100011001010011001001010100101100011001001111001010000; end
            14'd8438 : begin out <= 64'b1010001011010000101010100100110110100011010111010010100100011000; end
            14'd8439 : begin out <= 64'b1010010111111100101001100000011110011110101111011010001010001110; end
            14'd8440 : begin out <= 64'b1001110111001011101001100010111000011000110000111001101111011110; end
            14'd8441 : begin out <= 64'b0001111100010100001010101000011010101011011011010010010001110111; end
            14'd8442 : begin out <= 64'b1010100011001011101010111101111000100011101110111010001010111010; end
            14'd8443 : begin out <= 64'b0010101010000101000110100110100000100011001110001010100000101110; end
            14'd8444 : begin out <= 64'b1010101100000101001000010100110100100010110001011001111111100111; end
            14'd8445 : begin out <= 64'b0010101000101100000110010100101010011110001010111010001001011010; end
            14'd8446 : begin out <= 64'b0010001000001010101001001011100100101011011100100010011001011001; end
            14'd8447 : begin out <= 64'b1010001110001111001010101000011010101011100100000010100010001000; end
            14'd8448 : begin out <= 64'b0010010100000111001010111000000100100101101100001010100111101010; end
            14'd8449 : begin out <= 64'b1010000010011101001001101101000010100100111001110010101100100101; end
            14'd8450 : begin out <= 64'b1010100010110011001010100000011110101010001001011010100000001111; end
            14'd8451 : begin out <= 64'b0010101110110001101010110110000000101000011101100010100100000001; end
            14'd8452 : begin out <= 64'b1010000000101111101010001101101000001110100010001010101001111010; end
            14'd8453 : begin out <= 64'b1010011011011110001001000101010010101000011100100010011011001110; end
            14'd8454 : begin out <= 64'b1010000100100010101010101101101100101001110001011010011100001100; end
            14'd8455 : begin out <= 64'b0010100111000110001001010100101010100110111101110010101111010010; end
            14'd8456 : begin out <= 64'b1010011001010010001000000101111010101010111011001010100100110110; end
            14'd8457 : begin out <= 64'b1010001101000111101010100010001010100100000110111010010100100111; end
            14'd8458 : begin out <= 64'b0010010011100101001010110100111000100011111011111001110000111010; end
            14'd8459 : begin out <= 64'b1010101101110001101001011011000000100101101111011010101100100001; end
            14'd8460 : begin out <= 64'b0001010010110111101001110111110100100101101010010010011011000010; end
            14'd8461 : begin out <= 64'b1001110111001101101001100110001110101001011100010010100101001111; end
            14'd8462 : begin out <= 64'b0010000111100111001001100010100010100111101011001010100011001001; end
            14'd8463 : begin out <= 64'b0010100100000101001010110000101100011011111101011010011011110001; end
            14'd8464 : begin out <= 64'b1010011101011111001010111000001100101011101100111010100011110010; end
            14'd8465 : begin out <= 64'b1010011101111110001000110010100110100011001000111010101101001110; end
            14'd8466 : begin out <= 64'b0010100101101100101010111000000000101001110011011010101101101011; end
            14'd8467 : begin out <= 64'b1010011101100000001010100100011100100100011011101010011111001100; end
            14'd8468 : begin out <= 64'b1010101100111101001010101011100010101011101011011010100010010110; end
            14'd8469 : begin out <= 64'b0010101001100011101010100101101010101000111110101010101000010110; end
            14'd8470 : begin out <= 64'b0010011000100010001010111101010000011100110100001010100110011000; end
            14'd8471 : begin out <= 64'b0010001100100111001001110011101110100000100101100010010100100011; end
            14'd8472 : begin out <= 64'b0010010100110010001010000100111000101010100001101001110001111110; end
            14'd8473 : begin out <= 64'b0010000011111001101010111100010100100011010000101010101010010000; end
            14'd8474 : begin out <= 64'b0010101000101100101010011101111110100100010010101010011011110001; end
            14'd8475 : begin out <= 64'b1010100111100110101001110101111000101001110011111010100100000100; end
            14'd8476 : begin out <= 64'b0001110100101100001001101010110010101010111011100010010111001001; end
            14'd8477 : begin out <= 64'b1010100001110101101001000100111100100110111000000010101011100011; end
            14'd8478 : begin out <= 64'b1010101000001011001001010111100100100110110011010010101010111110; end
            14'd8479 : begin out <= 64'b0010101010111110001000010101001100011110110111111010101010110001; end
            14'd8480 : begin out <= 64'b0010011001000101100101101011101000101011111011010010011010110000; end
            14'd8481 : begin out <= 64'b1010100100000000001010011000000100101001011010000010010101100100; end
            14'd8482 : begin out <= 64'b1010010100011011101001001011110110101000111011110010101110111100; end
            14'd8483 : begin out <= 64'b0010101101111010001010001110000010101000100000001001011111010000; end
            14'd8484 : begin out <= 64'b0010011010101111100111101101100000100100001010110010010001110011; end
            14'd8485 : begin out <= 64'b1010110000000100101010100000001100010101011110011010001100101011; end
            14'd8486 : begin out <= 64'b1010001001010101101001110010000110101000100111111010001000110011; end
            14'd8487 : begin out <= 64'b0010100111001111001010011011000100101000011010011010100100110010; end
            14'd8488 : begin out <= 64'b0010100101101100101000011011000000101011100100010010100100111110; end
            14'd8489 : begin out <= 64'b1010010100001011101010100110110110101001110010100010011100111010; end
            14'd8490 : begin out <= 64'b0010101000000110001010011100011010101011011100001010100101010110; end
            14'd8491 : begin out <= 64'b0010010110000001000100011101011010100010010111000010010111010110; end
            14'd8492 : begin out <= 64'b1010101111101000101010101001011100100101001001101010011110101111; end
            14'd8493 : begin out <= 64'b1010101110000111101001010001100010011101100010001010100010001100; end
            14'd8494 : begin out <= 64'b0010000110111101001010111111100010101011011001010010101010001011; end
            14'd8495 : begin out <= 64'b1001110110111111001001001001001000101001110011010010010101010011; end
            14'd8496 : begin out <= 64'b1010100010110010001010011101100100100101010101011010101001010010; end
            14'd8497 : begin out <= 64'b0010011111011100001000110000000110101011011010011010101110100101; end
            14'd8498 : begin out <= 64'b0010101001100000101010100101110010100111110011011010010001010100; end
            14'd8499 : begin out <= 64'b0010101001001000101010011110110110100100110111100010010000010100; end
            14'd8500 : begin out <= 64'b0010101111001010101010010000011010011000101111111010101100101101; end
            14'd8501 : begin out <= 64'b1010010110111100001000010001011010010110110010001010101001100000; end
            14'd8502 : begin out <= 64'b0010010010011011100010100110011100101010011000011000001111011010; end
            14'd8503 : begin out <= 64'b0001110101011001001001100101001000100010101111001001110000111000; end
            14'd8504 : begin out <= 64'b0001110000101100001010100101011000101001100001010010110000001001; end
            14'd8505 : begin out <= 64'b1010100101011010001010111011111010101011101011101010001001110110; end
            14'd8506 : begin out <= 64'b1010100001000010100111111010000100101010110110010001100001110011; end
            14'd8507 : begin out <= 64'b0001111010111111001010001100010100101001110010100010100010110111; end
            14'd8508 : begin out <= 64'b0001111001100011001010111110110100100110010010100010101000011100; end
            14'd8509 : begin out <= 64'b0010010111101101101001010111001000010111011010100010101010101011; end
            14'd8510 : begin out <= 64'b1010100010010001001010110100010100100011111000111010101000001100; end
            14'd8511 : begin out <= 64'b1010101100110110101001001111000010100000111100000010010001100110; end
            14'd8512 : begin out <= 64'b0010100100011010001000000110100100101001000101000010100101101001; end
            14'd8513 : begin out <= 64'b1010000111001110101000100100011110101011110100111010101111100010; end
            14'd8514 : begin out <= 64'b1010101111000111101010010100010010101000101001000010100001111101; end
            14'd8515 : begin out <= 64'b1001010100110101101010100111111100101000011110101010001111010001; end
            14'd8516 : begin out <= 64'b1010101011110011001001100110010000100010001110110010100111110101; end
            14'd8517 : begin out <= 64'b0010100001100110101010101100000110100111001100111010010111100111; end
            14'd8518 : begin out <= 64'b0010000001010101000111000110101110100000011010010010001001110010; end
            14'd8519 : begin out <= 64'b0010011001010001001010101100111110101010001001001010010111011111; end
            14'd8520 : begin out <= 64'b1010010001110110001000001110001010100101111101001010011001011001; end
            14'd8521 : begin out <= 64'b0010010101110000101000011001110010101001110111101010101110101110; end
            14'd8522 : begin out <= 64'b0010010001001011001000001001011100101010110011111010101110011011; end
            14'd8523 : begin out <= 64'b1010000011100111001010011011010010101000001001001010101001111100; end
            14'd8524 : begin out <= 64'b1010100111111101101000011000001010100111110000010010011101100101; end
            14'd8525 : begin out <= 64'b0000111110010111001000010010001000011110100010010010101100110101; end
            14'd8526 : begin out <= 64'b1001111101111010101010111010011000101011011100100010100011111000; end
            14'd8527 : begin out <= 64'b1010101000101001101001001101000000100010101111110010110000001110; end
            14'd8528 : begin out <= 64'b1010010001010111101010101000111100101000110010011010000000100110; end
            14'd8529 : begin out <= 64'b1010101001000110101010001000010100100111001001010010001010010101; end
            14'd8530 : begin out <= 64'b1010100011011000001010010001110000101001111101011010101110101110; end
            14'd8531 : begin out <= 64'b0010000001111100101000011001010110101000001100000001011011010011; end
            14'd8532 : begin out <= 64'b1010010110101101001010001000100110011100100110101010000111010011; end
            14'd8533 : begin out <= 64'b0010100011100101101001111010100000100101011011110010100100000011; end
            14'd8534 : begin out <= 64'b1010011000111100101010011000100110100010111011100010101111000010; end
            14'd8535 : begin out <= 64'b0010101010111000101001010110010110101010100111000010101100110010; end
            14'd8536 : begin out <= 64'b0010010010010011101000000000001010100101011100101010100110111101; end
            14'd8537 : begin out <= 64'b0010010111010010001001011011001110100110111001000010010000100011; end
            14'd8538 : begin out <= 64'b0010110000000101000110110001111010100001011111110010100100011011; end
            14'd8539 : begin out <= 64'b1010001000110001001010101001111010101011111011111001000001101100; end
            14'd8540 : begin out <= 64'b1010010110101001101001001000011000101010001100100010000001000011; end
            14'd8541 : begin out <= 64'b1010000110100110001010111011111000101001011110101001111010100011; end
            14'd8542 : begin out <= 64'b0001011101101101101001110111000000100100011000110010100011010110; end
            14'd8543 : begin out <= 64'b0010101101111101001001111010110110100111110010011010101100010110; end
            14'd8544 : begin out <= 64'b0010101111111100101000011011010100101010010111110010100111100111; end
            14'd8545 : begin out <= 64'b0010101100100011001010111011111110100011010001111010000011100001; end
            14'd8546 : begin out <= 64'b1010101000100101001001101001000000101000100001010010011100101000; end
            14'd8547 : begin out <= 64'b0010001111111001101001010101110010101001010010101010100010011111; end
            14'd8548 : begin out <= 64'b1010010101111100101001011110010110100100110101100010101101011000; end
            14'd8549 : begin out <= 64'b1010011000111100101010111110111000101001111111100010101000111010; end
            14'd8550 : begin out <= 64'b1001111000110011000000000010111000101000011101101010001010101001; end
            14'd8551 : begin out <= 64'b1001101101110011001001110011001010101010101010100010011010000110; end
            14'd8552 : begin out <= 64'b0010101101100100001000101011001010100100011111010010100110111110; end
            14'd8553 : begin out <= 64'b1010101101000010101010011001101010101001000000110010000100101011; end
            14'd8554 : begin out <= 64'b0010101001010001001001100110101110101011000010000010001101101100; end
            14'd8555 : begin out <= 64'b1010101010101010101010111001010100100011001010001010100001000110; end
            14'd8556 : begin out <= 64'b1001010010111000101001010101100110101000011111100010100101101101; end
            14'd8557 : begin out <= 64'b0010100001110011100110101101001110101001110011011010100111001110; end
            14'd8558 : begin out <= 64'b0001110101101101100100011000100110101000111111111010110000001100; end
            14'd8559 : begin out <= 64'b0000101110010010001010011010111000101001011001111001111010000001; end
            14'd8560 : begin out <= 64'b0010011001110101000011010001100100101010011001111010100011101110; end
            14'd8561 : begin out <= 64'b1001110000111000001010011100000100101011101110110010010100000100; end
            14'd8562 : begin out <= 64'b1010100000010000100011100000010000101010010101011010011000111011; end
            14'd8563 : begin out <= 64'b0010100101001111001010111111101000100000110011101001110111011011; end
            14'd8564 : begin out <= 64'b1010101101010101101010100000010100101010001000000010100110000000; end
            14'd8565 : begin out <= 64'b0010101011100111001001010101011100101010010101010010100111001000; end
            14'd8566 : begin out <= 64'b1010100001010100001010010101111010101011111101111010101011110010; end
            14'd8567 : begin out <= 64'b0001100101001101001010110110100100101001111110001010100010000010; end
            14'd8568 : begin out <= 64'b1010010000110000101010101011101110101011000110001010101010101001; end
            14'd8569 : begin out <= 64'b0010101101000000101010001110010100101010010011100010101001010000; end
            14'd8570 : begin out <= 64'b0000010111001001101010010111110100100100011101111010011110010011; end
            14'd8571 : begin out <= 64'b1010100101110100001001001100101000101011100100110010101001000110; end
            14'd8572 : begin out <= 64'b1010011111000010001001001110110110101010110110010010100001110101; end
            14'd8573 : begin out <= 64'b1010100000110010001010010000000010101100000001100010011011101110; end
            14'd8574 : begin out <= 64'b0010010110000001001000101000100000101011111001100010011111001111; end
            14'd8575 : begin out <= 64'b0010000111000110101010100100010000101001111101001010101001101110; end
            14'd8576 : begin out <= 64'b0010011100100101001001101010011010101011100101110010000110100100; end
            14'd8577 : begin out <= 64'b1010101010001000001001010110100100101000001010011010010000101000; end
            14'd8578 : begin out <= 64'b0010101010000110101010001100110010100000100010010010100011110101; end
            14'd8579 : begin out <= 64'b0001111110110011001001011000100110101001001001101010101001010011; end
            14'd8580 : begin out <= 64'b0010010011000000001010101101001010100100101111100010011001011110; end
            14'd8581 : begin out <= 64'b1010100101011001001010100001011010101001100010001010010010000001; end
            14'd8582 : begin out <= 64'b0010101100111100101010010100101110101010110101000010110000100000; end
            14'd8583 : begin out <= 64'b1010101001011111001000100011101110101000110101100010011010111110; end
            14'd8584 : begin out <= 64'b1010101111001010101000100000010000100110011111011010010101000101; end
            14'd8585 : begin out <= 64'b0010100000100011101000100001000100100000111110110010101111000100; end
            14'd8586 : begin out <= 64'b0010000001000010101001011110101110101000010001001010100111001000; end
            14'd8587 : begin out <= 64'b0010100100100000001010011010110010101001010111011010100000110101; end
            14'd8588 : begin out <= 64'b0010010110100001101010001100100010100100001010011010100110001011; end
            14'd8589 : begin out <= 64'b1010001110101110001001101000001000100001001011100010001011011100; end
            14'd8590 : begin out <= 64'b1010010100001111001010011000010010100111001110101010101101001110; end
            14'd8591 : begin out <= 64'b1010100001001101001010100111100010011101111001100010011011101101; end
            14'd8592 : begin out <= 64'b0010101001010011101001101100001000100110001000110010101110001000; end
            14'd8593 : begin out <= 64'b0010101011111111101010111111010010100100101101011010101000101111; end
            14'd8594 : begin out <= 64'b0010001001010001001001111110110010100111011111011010101101011011; end
            14'd8595 : begin out <= 64'b1010100100101110101010011100001000100001000001110010100001000000; end
            14'd8596 : begin out <= 64'b1010010011110011001010010110011110101001100100001010011101100101; end
            14'd8597 : begin out <= 64'b0010010000101111101001000101011100100001111000110001100011010011; end
            14'd8598 : begin out <= 64'b1010101000101100101010101101010010100000000101001000001000101111; end
            14'd8599 : begin out <= 64'b1010100111101011101010110000000110101001111001110010100011111011; end
            14'd8600 : begin out <= 64'b0010101010001010001010101000101100101011000011110010100110011101; end
            14'd8601 : begin out <= 64'b0010010000111111001010110111001010100100100000110010010100011111; end
            14'd8602 : begin out <= 64'b0010101000100101001001101100111110101000001011010001101011011001; end
            14'd8603 : begin out <= 64'b0010101000011011001001000011000110100000100110110010101110101101; end
            14'd8604 : begin out <= 64'b0010000110101010001010111011010000101000111010011010011000111011; end
            14'd8605 : begin out <= 64'b0010011110011011001010100001111110100111011011000001101001011001; end
            14'd8606 : begin out <= 64'b0010101100110011101010011010100110101011010100100010001001001110; end
            14'd8607 : begin out <= 64'b0010101100001111001010110111100010011001001101111010101011011111; end
            14'd8608 : begin out <= 64'b1010100011001001001001110100111000101011101011000010011000101001; end
            14'd8609 : begin out <= 64'b0001110000101001101001110110100100100111010010011010101110100011; end
            14'd8610 : begin out <= 64'b0010101000111101001010010101111100101010101011111010101110010101; end
            14'd8611 : begin out <= 64'b1010101111001101100111110000111100101001100100001001101100111011; end
            14'd8612 : begin out <= 64'b0010100010001100001001101100000010101011000101110010101000101000; end
            14'd8613 : begin out <= 64'b0001110110011101101010111111101000011000100011001010101000101100; end
            14'd8614 : begin out <= 64'b0010100011011110100110101100001100010000010110011010010110101001; end
            14'd8615 : begin out <= 64'b0010010110000111001000010101111000011110010001110010101110001000; end
            14'd8616 : begin out <= 64'b1010011101011011101001100101101000101001101011010010101100011001; end
            14'd8617 : begin out <= 64'b0010101000111111101001001010110000101000111010101010100111110100; end
            14'd8618 : begin out <= 64'b0001100110011111001010000011000010100100011001100010100011011001; end
            14'd8619 : begin out <= 64'b0001010110000000001010101010001010100110010111001010010110100010; end
            14'd8620 : begin out <= 64'b0010010110001000101000010111110000101011001011011010000011111110; end
            14'd8621 : begin out <= 64'b1010011011010111101010000000010110100010101010000010100011100100; end
            14'd8622 : begin out <= 64'b0010100111101110001000001100000010100010000111010010101011111000; end
            14'd8623 : begin out <= 64'b1010101001010110101010111110011000100011011101010010100100110101; end
            14'd8624 : begin out <= 64'b0010011111000001101000100111000100100101101010001010011100000101; end
            14'd8625 : begin out <= 64'b0010101011110000000111001101100100011010101111001010100111111110; end
            14'd8626 : begin out <= 64'b0010000111001110101010101101011100011110110011101010100011101111; end
            14'd8627 : begin out <= 64'b1010010000101010101001011000000000100100111000001010101111001001; end
            14'd8628 : begin out <= 64'b1010101111111001001001101001001100101000001110101001110010110010; end
            14'd8629 : begin out <= 64'b0010101011110100001000000101001110100111101000110010101101010011; end
            14'd8630 : begin out <= 64'b1010011010000010000111011010000000101000010111110010010001011010; end
            14'd8631 : begin out <= 64'b0010100100100001101010000101100100101001001110010010010000000011; end
            14'd8632 : begin out <= 64'b0010010111000101000011110111001100100001101001111010101000011000; end
            14'd8633 : begin out <= 64'b1010001111010001001010100111000100100101001010001010100110111001; end
            14'd8634 : begin out <= 64'b0010011001101010001001110100011110100110101010000010001010011000; end
            14'd8635 : begin out <= 64'b0010010010011101101010111101010110100101101001111010100000110100; end
            14'd8636 : begin out <= 64'b1010000101101100001001010110011000100101111100001010101100000100; end
            14'd8637 : begin out <= 64'b0010100101011011101010000001111010101000010111010010000111001101; end
            14'd8638 : begin out <= 64'b0010100001001010001010110101111000100001000010110010010010101001; end
            14'd8639 : begin out <= 64'b1010100001101101000110100111001110010001101001011010100011110001; end
            14'd8640 : begin out <= 64'b0010010011001010101010010110000110100111010000001010010000100100; end
            14'd8641 : begin out <= 64'b1010001100110100100111101101111010101001101000001010100110100010; end
            14'd8642 : begin out <= 64'b0000100010110000001000011010110000101001101001101010010001110111; end
            14'd8643 : begin out <= 64'b1010100111001001000100110011110110101011011100000001100001110111; end
            14'd8644 : begin out <= 64'b1010001000101110001001111101111000100101011101000001011010110000; end
            14'd8645 : begin out <= 64'b1001000100100111001001100010011010100111110101110010011010010001; end
            14'd8646 : begin out <= 64'b0010100101010111101000000110111000100000011100001010010001010111; end
            14'd8647 : begin out <= 64'b0000110000110110101000001110100100101001001000011010100010110011; end
            14'd8648 : begin out <= 64'b1010101101001110001010110100001100101011111100001010100001010001; end
            14'd8649 : begin out <= 64'b0010010111001011001010000111010000101000101101000010011011000101; end
            14'd8650 : begin out <= 64'b0010100010110000101001000010100000101011110100000010010011101011; end
            14'd8651 : begin out <= 64'b1010010010000111000111101010010100100101100001011010011000010000; end
            14'd8652 : begin out <= 64'b0010010001010010101010001100000010100000000011000010011100011010; end
            14'd8653 : begin out <= 64'b1010101011001010101001000110010010101010110000110010100010110111; end
            14'd8654 : begin out <= 64'b0010001000011011001010100110010000101011101111010010010001110110; end
            14'd8655 : begin out <= 64'b0010000101000010001010111110000100100110001010010010001110001010; end
            14'd8656 : begin out <= 64'b1010100010100111100111011001111110100110111101010010001010111000; end
            14'd8657 : begin out <= 64'b0010011110011001100111001001011100100011111100000010100101111000; end
            14'd8658 : begin out <= 64'b1010101010101011101010000001111100101000010010101010100110110001; end
            14'd8659 : begin out <= 64'b1010100011100000101010110111111100011001010110111010100010100101; end
            14'd8660 : begin out <= 64'b0010100100100001001010010000110110011111100001010010001010110011; end
            14'd8661 : begin out <= 64'b1010101101010000101001011100110010101000010100110010001110011001; end
            14'd8662 : begin out <= 64'b1010101101011111001010101100100110100110000100110010010111110001; end
            14'd8663 : begin out <= 64'b0001111101001010101010001010111110101010101111000010101000001100; end
            14'd8664 : begin out <= 64'b1010000010001011001010010111110110100011001100011010011100111101; end
            14'd8665 : begin out <= 64'b1010010110000010101010111001100000100001110101011010010000111110; end
            14'd8666 : begin out <= 64'b0010101111100110001010100001100110001100101110111010101111101111; end
            14'd8667 : begin out <= 64'b1010010011111100101010011011101010100000101011100010101001101000; end
            14'd8668 : begin out <= 64'b1010011000101101001001001000000000101000110011001010101100010000; end
            14'd8669 : begin out <= 64'b1010011111011000101010100111011010101011110010100010100000101001; end
            14'd8670 : begin out <= 64'b0010001001001000101010100111101110100101011001011010010000101110; end
            14'd8671 : begin out <= 64'b1010100111000000001001100010010000101010111101101010101010111001; end
            14'd8672 : begin out <= 64'b0010101100101101101010000001000000100100010010101010100011101101; end
            14'd8673 : begin out <= 64'b0010011010111111001000101001110000101010010000011001110101011111; end
            14'd8674 : begin out <= 64'b1001111100000010101001111000010110100110110101001010101101011100; end
            14'd8675 : begin out <= 64'b1010010111001011101000011001010000100010011010000010000110101000; end
            14'd8676 : begin out <= 64'b1010011100111110101001010101000000101010001110110010101010010000; end
            14'd8677 : begin out <= 64'b1010101110000001101010000100110010101001011011110010100011100111; end
            14'd8678 : begin out <= 64'b0010001000001100001010010000010000100110111000011010001101001110; end
            14'd8679 : begin out <= 64'b0010011111011110000110101101001000100100101000010010100001010011; end
            14'd8680 : begin out <= 64'b1010101011011000000111101110011000100110111100011010100010101010; end
            14'd8681 : begin out <= 64'b1010010101001110101001111010101000101010001110101010100000110011; end
            14'd8682 : begin out <= 64'b1010001100101110101001110100010110101010110100110010101011001010; end
            14'd8683 : begin out <= 64'b1001111110110001101000000010100010101011001000100010100011010010; end
            14'd8684 : begin out <= 64'b1010101001111101001001110110001100101011001111110010101011101101; end
            14'd8685 : begin out <= 64'b1010101111101100101001011010111100011110101010100010011001010111; end
            14'd8686 : begin out <= 64'b0010100101001010101000001111111010101000101110000010100100000011; end
            14'd8687 : begin out <= 64'b0010101001111011001001110001010010101000010101011010100111110111; end
            14'd8688 : begin out <= 64'b1010100011110101001000111111110110101001010011011010011010100100; end
            14'd8689 : begin out <= 64'b0010100110101111001010101110011000100011001000011010100011000100; end
            14'd8690 : begin out <= 64'b1010101010000010001010001101000110101010101000001001101100001100; end
            14'd8691 : begin out <= 64'b0010100001111111001010000000110110100000111101100010100010110100; end
            14'd8692 : begin out <= 64'b1010000111001000001001101000001000100100001000011010101101011101; end
            14'd8693 : begin out <= 64'b0010000011110000001000111001100000101000101001111010101100010010; end
            14'd8694 : begin out <= 64'b0010000010001111101010100000101100100100010010000010100001111011; end
            14'd8695 : begin out <= 64'b1010101010001010101001000010000010011111011011111001110000110011; end
            14'd8696 : begin out <= 64'b0010100011111000000101000101000100010100011111010000111011000010; end
            14'd8697 : begin out <= 64'b1010101111001100101001011101001010100111001000101010010001011101; end
            14'd8698 : begin out <= 64'b0001110011010010101010011101111010010111001000011010001101110001; end
            14'd8699 : begin out <= 64'b1010000001110001001010111110101010100101110100111001100101110000; end
            14'd8700 : begin out <= 64'b1010101000000110101000111001000010101000010110111010101011011100; end
            14'd8701 : begin out <= 64'b1010100101110110001000000100000000101001101100010010011010001110; end
            14'd8702 : begin out <= 64'b0010101111110100101010110001100110010001111110010010100100111000; end
            14'd8703 : begin out <= 64'b0010001001010011001010110010010110101000101001110010100010110011; end
            14'd8704 : begin out <= 64'b0001111011100000001010011100001010101010111111100001110101011101; end
            14'd8705 : begin out <= 64'b0010101010001111001010001101010000100111000011110010000101101111; end
            14'd8706 : begin out <= 64'b1010011111100011001001101011111100101001010101110010010010111111; end
            14'd8707 : begin out <= 64'b0010100110100001100110110100001010101010100001000010000001110110; end
            14'd8708 : begin out <= 64'b1010100010110001001001100110100000100010011000011010000111010011; end
            14'd8709 : begin out <= 64'b0010100101111011001000110011101110101100001000100010011000010100; end
            14'd8710 : begin out <= 64'b1010100001111010001010101111000000101010101110100010100110001101; end
            14'd8711 : begin out <= 64'b0010010110111010001010010110011100100101010110011010101111001111; end
            14'd8712 : begin out <= 64'b0010101001000011001001100100110110101011000110110010011010010110; end
            14'd8713 : begin out <= 64'b0010001100011001001000011010010100100111111100101010101001000011; end
            14'd8714 : begin out <= 64'b0000110011001010001001110111111010100111100110100010010100000010; end
            14'd8715 : begin out <= 64'b1010010111101010001001011111100010101001110111001010101101001100; end
            14'd8716 : begin out <= 64'b1010010001111100101001010000010010101010101000101010100100111111; end
            14'd8717 : begin out <= 64'b1010101110100011001010011000100110101011010001101010011111111001; end
            14'd8718 : begin out <= 64'b0010000000011111001010001010110010101011111001110010100111111111; end
            14'd8719 : begin out <= 64'b1010010110110011001001100101110110100100000100100000110011011101; end
            14'd8720 : begin out <= 64'b1010101100111110101010100110101110100111100100100010100110111111; end
            14'd8721 : begin out <= 64'b1010010100110000001000010001110110101000010011101010100110011100; end
            14'd8722 : begin out <= 64'b0010001010110011100111011101010010101011001101010010101100111111; end
            14'd8723 : begin out <= 64'b0010010100101100001000011111011000101011000110010010100110101110; end
            14'd8724 : begin out <= 64'b0010011100111001101010010110011010101001100101000010010101100000; end
            14'd8725 : begin out <= 64'b0010101001100101001010001010111100101000001100010010011110100111; end
            14'd8726 : begin out <= 64'b1010010011111110001010000011101100100110100110011010100101000001; end
            14'd8727 : begin out <= 64'b1010101110001010101001100001011000100101000110011010101010110101; end
            14'd8728 : begin out <= 64'b0010100110010111101010100010111110101011101010100010010000101001; end
            14'd8729 : begin out <= 64'b0010100000101011101010011011100010101011111000110010010000111000; end
            14'd8730 : begin out <= 64'b1010100011001010100111111000010100101001101101010001110000000110; end
            14'd8731 : begin out <= 64'b0010011111001110101000010011110110101011101111010010011110000100; end
            14'd8732 : begin out <= 64'b0010100001101010001001001010010000100100100111101001101001000001; end
            14'd8733 : begin out <= 64'b1010011000110010001010001110010000100110100000010001111011110101; end
            14'd8734 : begin out <= 64'b1010100000111000101010110010110100101010001100001010100010111100; end
            14'd8735 : begin out <= 64'b0010010101100101101010110001010000100101110110111010101000111111; end
            14'd8736 : begin out <= 64'b0010100000011011101001101110111100101000101000010010011110100100; end
            14'd8737 : begin out <= 64'b0010101010010001101010010011110100100111100110110010100001010001; end
            14'd8738 : begin out <= 64'b0010011110011001001010000101111110101001011101010010001100000010; end
            14'd8739 : begin out <= 64'b1010010001100101101010001111000110101000000111010010010100010010; end
            14'd8740 : begin out <= 64'b1001110010010100101001110000111000101000010110110010101011111101; end
            14'd8741 : begin out <= 64'b1010101011010110101000010010111110101010001100010010011001100001; end
            14'd8742 : begin out <= 64'b0010010011011100001010101100010000101000100000010010100111000001; end
            14'd8743 : begin out <= 64'b0010011101101100001001011000110000101000111011101010101010110111; end
            14'd8744 : begin out <= 64'b1010010100101100001010100001110100100110001001110010000011101101; end
            14'd8745 : begin out <= 64'b0010100001000000101001001110000100101011111101100010101101010111; end
            14'd8746 : begin out <= 64'b1010011100100111101010000010111100100101011001010001110001011111; end
            14'd8747 : begin out <= 64'b0010001000010010001010000011101110101011110110001010101001011010; end
            14'd8748 : begin out <= 64'b0010101110011110001010110011001010100111101101010010011011010010; end
            14'd8749 : begin out <= 64'b1010011110001001101000111111110110101010101101000010100110111011; end
            14'd8750 : begin out <= 64'b1001111010111100101001001100001000101010101110011010101010000010; end
            14'd8751 : begin out <= 64'b0010100111010110101010101111010010100001010010000001111001111101; end
            14'd8752 : begin out <= 64'b0010100010101100101010010001011110011100011011010010100001110001; end
            14'd8753 : begin out <= 64'b1010100111000111001010100100100010101001010010010010100110001110; end
            14'd8754 : begin out <= 64'b0010011000010101101010101001111110100111010101111010100110101001; end
            14'd8755 : begin out <= 64'b0010101101111011001010100011010000100110101011110010011001011111; end
            14'd8756 : begin out <= 64'b1010011100111010001001101001101010100010111000110010100111110101; end
            14'd8757 : begin out <= 64'b1010010000110010001010011010110000101011101010111010101100000110; end
            14'd8758 : begin out <= 64'b0001101000000010001001100100111110101001101010010010011110101110; end
            14'd8759 : begin out <= 64'b0010101001110001001010101011001010011110110011100010101100100101; end
            14'd8760 : begin out <= 64'b0010100111101000101001100001001110100101100011001010011110101110; end
            14'd8761 : begin out <= 64'b0001110010101000001001100000100100101000110000001010100110011001; end
            14'd8762 : begin out <= 64'b0010101111111100001010001111110010100100000110111010100010010101; end
            14'd8763 : begin out <= 64'b0010100111101111101010101001000010101011010010010010010110101110; end
            14'd8764 : begin out <= 64'b1010011110000011101010110110010010100110011100101010100100000101; end
            14'd8765 : begin out <= 64'b1010101010111000101010001110000100010110011101000010001111010101; end
            14'd8766 : begin out <= 64'b0010000110000111101000111100001010100101001101001010101001100000; end
            14'd8767 : begin out <= 64'b0010101011101100101000110010011010101001101101101010000001011010; end
            14'd8768 : begin out <= 64'b0010011100111110101010101000000110011110110000000010010100110010; end
            14'd8769 : begin out <= 64'b0010101101010001001010110010001000101000001100001010011000101100; end
            14'd8770 : begin out <= 64'b0010100001100111101000100101111110100101000100000010100101001111; end
            14'd8771 : begin out <= 64'b1010001000100100001010100111011100100100101110111010000000101010; end
            14'd8772 : begin out <= 64'b0010101101110101001010000000000100011000100010111001111000101110; end
            14'd8773 : begin out <= 64'b0010101000110110001010010100010100000101010010111010101110000111; end
            14'd8774 : begin out <= 64'b0010100100001111101010100010010110101000110110101001100110001101; end
            14'd8775 : begin out <= 64'b0010100010100101001010011011010110101011001010101010100110011100; end
            14'd8776 : begin out <= 64'b0010010010010101001001100001010100101000110100001010011110101100; end
            14'd8777 : begin out <= 64'b0010100000111101101001111110010010101000101010100010010110001111; end
            14'd8778 : begin out <= 64'b0010011111010101001000000100011110101100010010001010011110000010; end
            14'd8779 : begin out <= 64'b1010010010101111100010000100101000100101000111111010110000000110; end
            14'd8780 : begin out <= 64'b0010100101010101001001010101101110101001000010001010011110110110; end
            14'd8781 : begin out <= 64'b0010011011000111001010011001111010011001101001111010100111100011; end
            14'd8782 : begin out <= 64'b1010101110111100001001000010001000100110001101111010010111001011; end
            14'd8783 : begin out <= 64'b0010100000000100101010001110011110100101110010110010011100000000; end
            14'd8784 : begin out <= 64'b0010000111001010101001111010000110101011110101000010010011100101; end
            14'd8785 : begin out <= 64'b0010010111111001101000010101111000100111001010101010100011101011; end
            14'd8786 : begin out <= 64'b0010000010011011001001011011111000101001001111101001111111111010; end
            14'd8787 : begin out <= 64'b1001111100110010101010111001011000101001100100011010001011011110; end
            14'd8788 : begin out <= 64'b0010010011100101001000010100011000100001001110010010100000101001; end
            14'd8789 : begin out <= 64'b1010101110110101001010100101010100101011101010000010011100000010; end
            14'd8790 : begin out <= 64'b1010010111111001001001110011011000101000100001010001100000011101; end
            14'd8791 : begin out <= 64'b1010101011010010001010101100100100100100101000101010010010101010; end
            14'd8792 : begin out <= 64'b1010101101010111101010011011011010101001000100001010010000111010; end
            14'd8793 : begin out <= 64'b1010101011100101000111011101010010011100100011010010010101001011; end
            14'd8794 : begin out <= 64'b1010101000011100101010100101111100010111001011000010000111111000; end
            14'd8795 : begin out <= 64'b1010101111100010101010000011111010101001101000110001110100110010; end
            14'd8796 : begin out <= 64'b1010001100001100001010000010011100100110000110000001111101001010; end
            14'd8797 : begin out <= 64'b0010010101011110101010010000101000011100111010101010101111100010; end
            14'd8798 : begin out <= 64'b1010100111101001001010101010101000101001001101010010011000110000; end
            14'd8799 : begin out <= 64'b1010011110001101101010101100111100100111010101010010000010001011; end
            14'd8800 : begin out <= 64'b0010101101000010001001000111110000100110101101101001101010000111; end
            14'd8801 : begin out <= 64'b1001010001001111101010101000010000101001100110111010010101101110; end
            14'd8802 : begin out <= 64'b0001111110010110101010100101001110101011010001101010101011001000; end
            14'd8803 : begin out <= 64'b0010101001010010001001001111100100010101011111010010101111000111; end
            14'd8804 : begin out <= 64'b1001011001101101001010010001110010100111111111101010101101101010; end
            14'd8805 : begin out <= 64'b0010101100111110101010100000010000011000010100001010011001000100; end
            14'd8806 : begin out <= 64'b0001111101101000001010100100001000101000001111011010100010000011; end
            14'd8807 : begin out <= 64'b1010101011001100101001010000110000100110011100101010000001010111; end
            14'd8808 : begin out <= 64'b0010101010101000101010001100101010100001101101001001110100100101; end
            14'd8809 : begin out <= 64'b1010100000101011001010011111101100101100001101101010101101110000; end
            14'd8810 : begin out <= 64'b0010100100001001101010011101100110101011000111010010101010010101; end
            14'd8811 : begin out <= 64'b0010101101110100101010100100011100101001101000001010101101110110; end
            14'd8812 : begin out <= 64'b0010001101110011101001010001110010101000011101100010100001101001; end
            14'd8813 : begin out <= 64'b0010100000000000101010001110011000101000011010110010011011011110; end
            14'd8814 : begin out <= 64'b0010100101100100101001010111000100100101000100111010101111001010; end
            14'd8815 : begin out <= 64'b1010100011101100001001100101011010101010111001101010010001110011; end
            14'd8816 : begin out <= 64'b0010011011000010001010100010011110100101000101010010100001110110; end
            14'd8817 : begin out <= 64'b1010101010101000001001101000001100100110100111100010101001111111; end
            14'd8818 : begin out <= 64'b1010101100100110001010101101101000011101000011001010011100111110; end
            14'd8819 : begin out <= 64'b1010101011010100101010110011000100101001100100101010011111000011; end
            14'd8820 : begin out <= 64'b0010010100101111101010010111010100100010010111110010100001010010; end
            14'd8821 : begin out <= 64'b0010101111110000000111010011111000100100001110101010101010001111; end
            14'd8822 : begin out <= 64'b1010100101100011001001001111100110011101011110010010101011101011; end
            14'd8823 : begin out <= 64'b1010001110100110001000100011111110100101110010100010010100110110; end
            14'd8824 : begin out <= 64'b0010101100111101100110000110001010101011110011011010101011101110; end
            14'd8825 : begin out <= 64'b1000010111101101101010011000010110101100000100111001110011110010; end
            14'd8826 : begin out <= 64'b1010101000010011101001000000101010011101001101111010101000001011; end
            14'd8827 : begin out <= 64'b1010101000110011101000110101111000101011101101100010101000010001; end
            14'd8828 : begin out <= 64'b1010011000101010000111100010011100101011110111001010101110000010; end
            14'd8829 : begin out <= 64'b0010010110101101000100111011100010100100001000000010100000101001; end
            14'd8830 : begin out <= 64'b1010100101010011001010001100100100101001101000010001111000001011; end
            14'd8831 : begin out <= 64'b1010001010001001000111000111001010100010111100110010100101000110; end
            14'd8832 : begin out <= 64'b1010000110010000101010110000001100101010011111001010100110100001; end
            14'd8833 : begin out <= 64'b0010101011100110001001110001001000101011010101011010100001011110; end
            14'd8834 : begin out <= 64'b1010010100000110001010110010110110100001111011111000010100011001; end
            14'd8835 : begin out <= 64'b0010100100100011101010100010101100100111001010001010010000001000; end
            14'd8836 : begin out <= 64'b0010100001010000100111000010011110101001000111111010011000001011; end
            14'd8837 : begin out <= 64'b1010100010011001101010010000100110100100111100011001011110100001; end
            14'd8838 : begin out <= 64'b1010011101001000001010100010100000100100111011001010100001110111; end
            14'd8839 : begin out <= 64'b0010100001101000101001000001010110101000000010010010101011100110; end
            14'd8840 : begin out <= 64'b1010011111000101100110110011010110001110111110000010100011011010; end
            14'd8841 : begin out <= 64'b1010000010010011001001011010101100100110101001011001001110000000; end
            14'd8842 : begin out <= 64'b1001111111110101101000101011110100101011111110000010010001101000; end
            14'd8843 : begin out <= 64'b0001011011001110001010001111101100100100000001100010010011000110; end
            14'd8844 : begin out <= 64'b0010100101100001001010100100100000101010000101101010100000010001; end
            14'd8845 : begin out <= 64'b0010011111101001001010001100101100100001000101011010100110110001; end
            14'd8846 : begin out <= 64'b1010100001110100101001010110110010100100101101010010010011000000; end
            14'd8847 : begin out <= 64'b0010100110000101001010110101001100100110001000000010100011110000; end
            14'd8848 : begin out <= 64'b1010100111010010100110101010110010101001010010100001100101010001; end
            14'd8849 : begin out <= 64'b1010100111111010001010111101011000101010111111101010101100100011; end
            14'd8850 : begin out <= 64'b0001001011111000100111111100100110101011100010000010011100100001; end
            14'd8851 : begin out <= 64'b0010011111100001001000111011000000101000101011001010011000100000; end
            14'd8852 : begin out <= 64'b1010011000010000001001110110111100100100011101110010110000000011; end
            14'd8853 : begin out <= 64'b0001111100111111001010001010101000100010011100001001111001101111; end
            14'd8854 : begin out <= 64'b1010010000100001101001010000111000011100000101011010000110101010; end
            14'd8855 : begin out <= 64'b0010001111010111001010000011010010101011111011011010011001011101; end
            14'd8856 : begin out <= 64'b1010000101011100101010100111101010101001110101001010011100000111; end
            14'd8857 : begin out <= 64'b1010100111011101001010111111000110100010101100000010101010010101; end
            14'd8858 : begin out <= 64'b0001111010111010101010001111001100100101011101011010011010000111; end
            14'd8859 : begin out <= 64'b1010010101010111001010101101001110101000000100010010011101010100; end
            14'd8860 : begin out <= 64'b0010101011110011101001110110101000011001001010110010010001001100; end
            14'd8861 : begin out <= 64'b0010010110111010001001110111010000100110110001010001001000110010; end
            14'd8862 : begin out <= 64'b1010000101001110001000100101101000011110010100110010101010000110; end
            14'd8863 : begin out <= 64'b1010001110110110101000000000010000101001010001000010101000011100; end
            14'd8864 : begin out <= 64'b0010101000001000101010100000111000101011101111111010010110110101; end
            14'd8865 : begin out <= 64'b0001000100100100101010100001100100101011000001010010100111101001; end
            14'd8866 : begin out <= 64'b1010010000011111001010010111010010101000100000101010101100000010; end
            14'd8867 : begin out <= 64'b0010100101100000001000010011000000101011101110001001011011101010; end
            14'd8868 : begin out <= 64'b1010100100000111101010001000011110011111000110010010101010011000; end
            14'd8869 : begin out <= 64'b0010011000101010101010010011111010101010000011101010100000001011; end
            14'd8870 : begin out <= 64'b0010011111110011001010100111101100101000000111001010100001010000; end
            14'd8871 : begin out <= 64'b0010010010100110001001000010101010100111000010001010101010001111; end
            14'd8872 : begin out <= 64'b0010101101001011001010100001101100011010100101101010010101000101; end
            14'd8873 : begin out <= 64'b0010101000000000001010011010010010101000000001010010001101111110; end
            14'd8874 : begin out <= 64'b1010010011111111101010011101001000101001101010001010010100111001; end
            14'd8875 : begin out <= 64'b0010100011011100101001111010010010100110011001001010100011001001; end
            14'd8876 : begin out <= 64'b0010100011010100001001110100011110101001011110011010110000010110; end
            14'd8877 : begin out <= 64'b1010100110101110101000101001000010100111100110111010010111100001; end
            14'd8878 : begin out <= 64'b0010001110000011100111001110000000101010110001100001100110011100; end
            14'd8879 : begin out <= 64'b0001111101000110101010011001001000100101010110001010101001111110; end
            14'd8880 : begin out <= 64'b0010011010001111100110000010000000101011110111101010010100100110; end
            14'd8881 : begin out <= 64'b1010100101100111101010111010110100101010000101110001100010001111; end
            14'd8882 : begin out <= 64'b1001110000101001001010000110010000101011100011110010100000000101; end
            14'd8883 : begin out <= 64'b1010100111100011001010000110000100101010011111010010100111101100; end
            14'd8884 : begin out <= 64'b1001100101101111001010100000111000011000111110110010101101110101; end
            14'd8885 : begin out <= 64'b0001111010000001101001100110000100100111000101100010101001011101; end
            14'd8886 : begin out <= 64'b1010010101000011001001100101110100101001110110001010101010110101; end
            14'd8887 : begin out <= 64'b1010011111010011101001110000010110100011111110110001111111110101; end
            14'd8888 : begin out <= 64'b0010011010101101001001110101100000011110010111011010000110001000; end
            14'd8889 : begin out <= 64'b1010101000110111001010010000100010101001110110001010101011001111; end
            14'd8890 : begin out <= 64'b1010101011101110101010000111101010100110110011010010101100101001; end
            14'd8891 : begin out <= 64'b1010010001001100101010110100010000101010000000001010101101001011; end
            14'd8892 : begin out <= 64'b0010100110000000001000110100100010011101011101010010101100101100; end
            14'd8893 : begin out <= 64'b1010010011100001101010011011100110100011001001000010001101011000; end
            14'd8894 : begin out <= 64'b0010101000010111101010011101001110100000111100000010100100110110; end
            14'd8895 : begin out <= 64'b0010101100010110101010010010101010100011100001111010010111010001; end
            14'd8896 : begin out <= 64'b0010101000011001101000010111010110100000110111100001110101010010; end
            14'd8897 : begin out <= 64'b1010100100010110000110101111111000101011010100100010000100100110; end
            14'd8898 : begin out <= 64'b0010100100000001101001010101101100011101111111011010001111110111; end
            14'd8899 : begin out <= 64'b1010100100011101101010111010000010101010110100111010011111010000; end
            14'd8900 : begin out <= 64'b1010101110100010101001001001100010100110000011100010010001001000; end
            14'd8901 : begin out <= 64'b0010001100101101001001110100001100100101111000100010010101100010; end
            14'd8902 : begin out <= 64'b0010001010101100001000111000101100101000010011001010011010000110; end
            14'd8903 : begin out <= 64'b0010011111100010001001011011100010101000110000110010000101110000; end
            14'd8904 : begin out <= 64'b1010010111100101001010010000001000010111010010010010100001100010; end
            14'd8905 : begin out <= 64'b1010100011100001100111110001101010100010101011001010100111010111; end
            14'd8906 : begin out <= 64'b0010101000011011001010010000100010101000100000110010101110000011; end
            14'd8907 : begin out <= 64'b0010100001110001001010101010101110100010010001011010010111011100; end
            14'd8908 : begin out <= 64'b1010101110100101001000001101011100011110001000111010010000101000; end
            14'd8909 : begin out <= 64'b0001110100001001101010001001001110100101011011011010000110110111; end
            14'd8910 : begin out <= 64'b1010011110001101101010101001000100101010001101101001100010110100; end
            14'd8911 : begin out <= 64'b0010010111100000101010001010011000100011000101110001111110111001; end
            14'd8912 : begin out <= 64'b1010101100011110101000111100101110100001011110111010101100111111; end
            14'd8913 : begin out <= 64'b1001111110011001101001111100011110101000001101000010000100010100; end
            14'd8914 : begin out <= 64'b0010000110100001001001100011111000101011001000001010010011100001; end
            14'd8915 : begin out <= 64'b1001100101100111001001100011010010011101111111101010101001000100; end
            14'd8916 : begin out <= 64'b0010100100111100000110101010100100001100011001101010101110011100; end
            14'd8917 : begin out <= 64'b0010101110100111101010111110011000100100111010101010101101011000; end
            14'd8918 : begin out <= 64'b0010011101101011101010010011011100100101001010100010011101000111; end
            14'd8919 : begin out <= 64'b0010101111010101001000000111111000101001010011111001000100010100; end
            14'd8920 : begin out <= 64'b0010101011000011100111001110001000100010100101100010101001011110; end
            14'd8921 : begin out <= 64'b0010010011111000001010101010110100101100000101011001010010111000; end
            14'd8922 : begin out <= 64'b1010100110100111101010001101000110011000011101001010000111011100; end
            14'd8923 : begin out <= 64'b0010101111010010001010011101000100100000010001010001110110100010; end
            14'd8924 : begin out <= 64'b1010100110011010001010111001110100100111001000010010011101110100; end
            14'd8925 : begin out <= 64'b1010101001000001101010011001010010101000101110100010001001010101; end
            14'd8926 : begin out <= 64'b1010101110111011101001011010001110101001010101011010101110111000; end
            14'd8927 : begin out <= 64'b0010101100111001001010110011001010101001010101011010100010100011; end
            14'd8928 : begin out <= 64'b0010100110010110101010110101010100100001011001110010100000000001; end
            14'd8929 : begin out <= 64'b0010100000111011000110111110011010101011101000001010010111100011; end
            14'd8930 : begin out <= 64'b1010000100000110100110000100111110011101010111001010001001000110; end
            14'd8931 : begin out <= 64'b0010101000001010001000011111001100100100101000001010011100111110; end
            14'd8932 : begin out <= 64'b0010101001110001001010011000101010100000101111101010100010000101; end
            14'd8933 : begin out <= 64'b1010100101110010101010100111001000011101110110110010000101100110; end
            14'd8934 : begin out <= 64'b1010101000000000101010000000010000101001011101011010101111101110; end
            14'd8935 : begin out <= 64'b1010010011000001101010000101111000000000100100110010100010101011; end
            14'd8936 : begin out <= 64'b0010101000011011001000111110000010100110101000101010100010100000; end
            14'd8937 : begin out <= 64'b0010011000011000001000010101100000011101000001100010100101011001; end
            14'd8938 : begin out <= 64'b0010000001000010001001010111001100101011000000101010011100111101; end
            14'd8939 : begin out <= 64'b1010011001010011001000111111111010101011011111100010010111111000; end
            14'd8940 : begin out <= 64'b0010011011000000101010111101110000101100000100101010100111100001; end
            14'd8941 : begin out <= 64'b0010010010111111001000110010100110101011110010110010101001001110; end
            14'd8942 : begin out <= 64'b1010101101100111001001001011101100101010110101000001111101100110; end
            14'd8943 : begin out <= 64'b0001010000101001001010111101000100101010101100010010010001100010; end
            14'd8944 : begin out <= 64'b1010011110010010001010111101100100101010110110000001110001001000; end
            14'd8945 : begin out <= 64'b0001111000100000100110100011100000101011101101111010011000011100; end
            14'd8946 : begin out <= 64'b0010011010100001001001001111010010100000110010011010010110001110; end
            14'd8947 : begin out <= 64'b0010101001110100001000001000101010100001001110111001111100111100; end
            14'd8948 : begin out <= 64'b1010100100011001100111110000011010100101001011011010100111101100; end
            14'd8949 : begin out <= 64'b0010100001010000001010000101011000101001100100010010101110001001; end
            14'd8950 : begin out <= 64'b0010010100110010101010000111011010101000010001111010101000010010; end
            14'd8951 : begin out <= 64'b1010000000100001101010010110110100100101010110010010101101101011; end
            14'd8952 : begin out <= 64'b1010100000001011101010111111001100100111010000101010101101010110; end
            14'd8953 : begin out <= 64'b1010010000110110001010101010001010100001001001011010101001010101; end
            14'd8954 : begin out <= 64'b0010100101111001101010000010001100100101010000101001111000111000; end
            14'd8955 : begin out <= 64'b0010011100001111101001101110011110101000000001110010100100010101; end
            14'd8956 : begin out <= 64'b1010100011110001101001111000001110100110000110011010101101110100; end
            14'd8957 : begin out <= 64'b1010100100100100101010100000100100100101110011101001110010111011; end
            14'd8958 : begin out <= 64'b0010101100101010001010110111100000100101111101111010011000011000; end
            14'd8959 : begin out <= 64'b0010101000111010101010101110010010100010100101001001111100100100; end
            14'd8960 : begin out <= 64'b1010100001010010001001000110101010100010000010111010100110011000; end
            14'd8961 : begin out <= 64'b0010100010101110101001111111010110101001111110000001010100100110; end
            14'd8962 : begin out <= 64'b0010101011101101000111110011111000101001111100010010100010111000; end
            14'd8963 : begin out <= 64'b0010101001011111001011000001011010100010111001101010000010011010; end
            14'd8964 : begin out <= 64'b0010011000111010001001100010011110101000101111110010101000101001; end
            14'd8965 : begin out <= 64'b1010100100011100000111111100001110101001001001100010100110100010; end
            14'd8966 : begin out <= 64'b1010101100110000001010111111001110100100010101011010010101101110; end
            14'd8967 : begin out <= 64'b1010010101110010101010101101111000101001010110010010101111001110; end
            14'd8968 : begin out <= 64'b0010011100011101001001000111010010100010000001010010100011001000; end
            14'd8969 : begin out <= 64'b0010001111011100100010001001001000100001100011100010100101011011; end
            14'd8970 : begin out <= 64'b0010101110000111001010001100100000101011000110010010101111000011; end
            14'd8971 : begin out <= 64'b1010101110111010101010001100111000101001001000010010010110011110; end
            14'd8972 : begin out <= 64'b0010001111110110001010000110110110101000011111100001100000011100; end
            14'd8973 : begin out <= 64'b1010100010011101101010101100100010101001010001111010100111111110; end
            14'd8974 : begin out <= 64'b0010100001011110001001001100101010101000110001000010101110000100; end
            14'd8975 : begin out <= 64'b1010010110111101001000101000010110100111110000001010010001010000; end
            14'd8976 : begin out <= 64'b0010010010111010101010000010001100101001101111000010000110111010; end
            14'd8977 : begin out <= 64'b1001110111100000101001001100000110100100111110010010101101110010; end
            14'd8978 : begin out <= 64'b1010100011000010001001111010000010101011111111100010101110000010; end
            14'd8979 : begin out <= 64'b0010100010111011101010100110010110100110001001100010101010110100; end
            14'd8980 : begin out <= 64'b1010100010010111101001100011101010100011011011111001110011100101; end
            14'd8981 : begin out <= 64'b1010000011001000001001011000111010011110010010000010100011110110; end
            14'd8982 : begin out <= 64'b0010000100001110001010011001011010100110101101011001101100101000; end
            14'd8983 : begin out <= 64'b0001111110111011101010010010001110100110101010110010010011100110; end
            14'd8984 : begin out <= 64'b0010010111100101100111100110010100011111010110000010011101110101; end
            14'd8985 : begin out <= 64'b0010000110001101100110101010010100100111101010111010101100001010; end
            14'd8986 : begin out <= 64'b0010010110100000100110101101000100101100000011011010011110001001; end
            14'd8987 : begin out <= 64'b1010100100110001000100001011000100100100000001100010011010000001; end
            14'd8988 : begin out <= 64'b0010000100000010101001010110000100100000010000010001110101100111; end
            14'd8989 : begin out <= 64'b0010010111101111001001101100011000100101010001001010011110100010; end
            14'd8990 : begin out <= 64'b0001110010001000001011000010111100101001000111100010100001000110; end
            14'd8991 : begin out <= 64'b1010101101010000101001010101110110100110100000011001100100101010; end
            14'd8992 : begin out <= 64'b0010011001111010101001101100011010101001000111010010000110111100; end
            14'd8993 : begin out <= 64'b0010101000000010101000111101011100100100111101111010101100101011; end
            14'd8994 : begin out <= 64'b1010101110010100001000000011101100101010110011000010100011100101; end
            14'd8995 : begin out <= 64'b0010100011100011001010001010011110100000001010010010100011010110; end
            14'd8996 : begin out <= 64'b0001111100000001001010011001101010001110001111100010011010011001; end
            14'd8997 : begin out <= 64'b0010011111000010001000000100010100101010011100111010100000110100; end
            14'd8998 : begin out <= 64'b0010101110101001101010110011000000101000100010001010010101100011; end
            14'd8999 : begin out <= 64'b1010100010001011001010101110001110100010110010111010011110001111; end
            14'd9000 : begin out <= 64'b0010101101100000001000000110110010100011001100001010101011000010; end
            14'd9001 : begin out <= 64'b1010101010100111101010111101001000101000000000111010101101101001; end
            14'd9002 : begin out <= 64'b1001111110011000101000111111000100100000011100111010100111001101; end
            14'd9003 : begin out <= 64'b0010100110100011001001110000110110100011010110100010101101110111; end
            14'd9004 : begin out <= 64'b0010101110011000101001101111001100100110011001000010010000110100; end
            14'd9005 : begin out <= 64'b1010010000001111101001010000110100101011010010001010011110011010; end
            14'd9006 : begin out <= 64'b0010100100110111001001110011111100101010100110000010010001000000; end
            14'd9007 : begin out <= 64'b0010100111011100001011000011011100100010111100100010100000110111; end
            14'd9008 : begin out <= 64'b1010101111111011101010010110100100011111010011010010000110111010; end
            14'd9009 : begin out <= 64'b1010100011001101001000001001100110101010001010010010100111001001; end
            14'd9010 : begin out <= 64'b0001111000011101001001110010110110101011000101010010101111100101; end
            14'd9011 : begin out <= 64'b0010011000101011000111010111000100011100100010110010010101011111; end
            14'd9012 : begin out <= 64'b0010011110011111101000110101110110011110110111101010011011110000; end
            14'd9013 : begin out <= 64'b0010100011001001101001101001111110100100001010111010100011100010; end
            14'd9014 : begin out <= 64'b0010011000000010100101111010011110100110001011100010100001101110; end
            14'd9015 : begin out <= 64'b0010001001101111101000111010111010100010110001111010100111111001; end
            14'd9016 : begin out <= 64'b0001001000010010001010101011011100101011110110110010100111110011; end
            14'd9017 : begin out <= 64'b0010100110110111000111111111111010101010010001110001100001101001; end
            14'd9018 : begin out <= 64'b1010011010001000101010111001100110101010101001010001111001110100; end
            14'd9019 : begin out <= 64'b1010001100001110001010001110011110101000000001100001011011010001; end
            14'd9020 : begin out <= 64'b0010011010010111001010001011111000100110000110010010101001011011; end
            14'd9021 : begin out <= 64'b0010100011000001000111010110011000100001011110001010101100100010; end
            14'd9022 : begin out <= 64'b0010100011111001101010001010110000101000111011101010101110011010; end
            14'd9023 : begin out <= 64'b0001001001011110001010000101000000101001111111101010001111111010; end
            14'd9024 : begin out <= 64'b0010011100110000101001010000000110011100001111001010101110010101; end
            14'd9025 : begin out <= 64'b1010101001111011101010100011100010011000011001110010100101101110; end
            14'd9026 : begin out <= 64'b1001110110111111001001011001010100101011100011010010010100001010; end
            14'd9027 : begin out <= 64'b0010100001001100101010011001001110100110001101011010100110001111; end
            14'd9028 : begin out <= 64'b0010101000111011001010011101010010101001111100001010101111011001; end
            14'd9029 : begin out <= 64'b0010000110101010001010110111010100100110000011001010101011000100; end
            14'd9030 : begin out <= 64'b0001111001011001101000011110001110100111110001110010100000100001; end
            14'd9031 : begin out <= 64'b0010010110101010100111111111111110101000011000010010010001011101; end
            14'd9032 : begin out <= 64'b0010010011100100001001100101010000101000010000011010011100100111; end
            14'd9033 : begin out <= 64'b0010100100110110001001011011011000101010111110000010000100000000; end
            14'd9034 : begin out <= 64'b0010011100000111001010001001111110101000000011000010001011011001; end
            14'd9035 : begin out <= 64'b1010011010110000101010000101001100101000111110101010100011100000; end
            14'd9036 : begin out <= 64'b0010100011100101101001011001101000101000001001011010100110011001; end
            14'd9037 : begin out <= 64'b0010100100111001101000011000110010101001011101011010100011111111; end
            14'd9038 : begin out <= 64'b1010101111011111001010100010010010100100101101110010100000011100; end
            14'd9039 : begin out <= 64'b0010101100101110001010100111110010010000110010000010010110010110; end
            14'd9040 : begin out <= 64'b0010100010001011100111110100011000101011111011001010100100100111; end
            14'd9041 : begin out <= 64'b1001111111101010101010101100101100100000100100111010100100101111; end
            14'd9042 : begin out <= 64'b1010100100011011100111001101011100100101111110011010100011100110; end
            14'd9043 : begin out <= 64'b1010011000100110100110000000101000101010000110000010101010010101; end
            14'd9044 : begin out <= 64'b1010100010101100001010111001100110101000100110110010101000111101; end
            14'd9045 : begin out <= 64'b0010011011011100001010000111111110101011101110011010101000001000; end
            14'd9046 : begin out <= 64'b1010010010010100001010010100111000101010111001011010010100110110; end
            14'd9047 : begin out <= 64'b1010010011101000101001001000011010101000001001111010100000011001; end
            14'd9048 : begin out <= 64'b1010100111010001001001101100010100101010111100010010101111101100; end
            14'd9049 : begin out <= 64'b0010010000101011101001111110100100100110110100010010011100111001; end
            14'd9050 : begin out <= 64'b1010011101101110101010111001001100100110101000001010010001111001; end
            14'd9051 : begin out <= 64'b0010101000100010001010111101101110101001000000100010011100110100; end
            14'd9052 : begin out <= 64'b1010010011101101001001000111101100010111110101010010101110010010; end
            14'd9053 : begin out <= 64'b0010010110000010101010001010011110100010000111001010100010101011; end
            14'd9054 : begin out <= 64'b0010101011100000101010000110111110011110011110111010100110110011; end
            14'd9055 : begin out <= 64'b1010000100101101001010011011010000101011001101011010101101000001; end
            14'd9056 : begin out <= 64'b0010100111010000101000001001011010100101000010100010010100111100; end
            14'd9057 : begin out <= 64'b1010101011100111101000100001111000100110110101101010101111100011; end
            14'd9058 : begin out <= 64'b0010101101011011101001001001011010101010010111011010101011000100; end
            14'd9059 : begin out <= 64'b1001111000110110001010101111011100101010101110100010101010101011; end
            14'd9060 : begin out <= 64'b1001100011111000001010111011001110101001110101000010100011010111; end
            14'd9061 : begin out <= 64'b0010010010001010100110110111010110100100110100101010101011100000; end
            14'd9062 : begin out <= 64'b1010101100011010100111000111010000100111111000110010010011000000; end
            14'd9063 : begin out <= 64'b0010101101000001101010001110011000100000010100001010010101001110; end
            14'd9064 : begin out <= 64'b1010100010100100101011000101000010100100100101000010011010011011; end
            14'd9065 : begin out <= 64'b1010010111000110001010111110111000100010110110001010011011000011; end
            14'd9066 : begin out <= 64'b1010010001001101001001100101000110101000000011100010101011101110; end
            14'd9067 : begin out <= 64'b1010101000101110001001101111010010100110100111000010100110001000; end
            14'd9068 : begin out <= 64'b1010100001011010001000000111000100101000010100101010100100011110; end
            14'd9069 : begin out <= 64'b1010101010100100101001110101100000101010111000110010010000000110; end
            14'd9070 : begin out <= 64'b1010100011000110101010101001001110101010111110000010100111011100; end
            14'd9071 : begin out <= 64'b0010011110110110101010110101110110100111001110011010011001100100; end
            14'd9072 : begin out <= 64'b1001101001011101101010100001111100100001110110110010100101101000; end
            14'd9073 : begin out <= 64'b1010101110010010101001101010001100100011011010111010010101000111; end
            14'd9074 : begin out <= 64'b1010001001010010101000011011010110100110000010000010101000111101; end
            14'd9075 : begin out <= 64'b0010100111110110001000111100000110100100101001100010100010111010; end
            14'd9076 : begin out <= 64'b1010101001011010000111100001000110100111000001000010101101101110; end
            14'd9077 : begin out <= 64'b0010100101001111001010001101010100100110011111001010100100110110; end
            14'd9078 : begin out <= 64'b0010011010110101101010011000011110101001110000110010010100111100; end
            14'd9079 : begin out <= 64'b1010001000011111001001100011100000101001111001001001111000000010; end
            14'd9080 : begin out <= 64'b1010101101001101101010100001011010011001010011001010010100111111; end
            14'd9081 : begin out <= 64'b1010011001100000001001110110101110011001011101110010100010000011; end
            14'd9082 : begin out <= 64'b0001110101101110001001001010001000101011010010000010001111100100; end
            14'd9083 : begin out <= 64'b0010000001101011001010000010110010100101000111010010010011101001; end
            14'd9084 : begin out <= 64'b1000000101110110001000010000011100100111101000000010101010111011; end
            14'd9085 : begin out <= 64'b1010101111000010001000100100101100010110010101111010001001011101; end
            14'd9086 : begin out <= 64'b1010101001011011001001110110000100100101001101100010100000001111; end
            14'd9087 : begin out <= 64'b0010101100110011101001001010001000100111000000000010010101110000; end
            14'd9088 : begin out <= 64'b0010100000010010001011000010000110101001100011111010101111010000; end
            14'd9089 : begin out <= 64'b1010000001001110001010111001001110100100001100011010011101101101; end
            14'd9090 : begin out <= 64'b0010001001011010001010001011000000100100001111110010101011100110; end
            14'd9091 : begin out <= 64'b0010100000110100001010111101110000011111010011111010001101011001; end
            14'd9092 : begin out <= 64'b1010010000000000101001000010100100101000111001011010100111010000; end
            14'd9093 : begin out <= 64'b1010101011110010100110011101100010101010010011111010101110100110; end
            14'd9094 : begin out <= 64'b1001100110000111001010101110111000100101111101010010100000111011; end
            14'd9095 : begin out <= 64'b0010010000110010100101100001110110101011100110010010100001010001; end
            14'd9096 : begin out <= 64'b1010100110101111001001010011111010100100000110100010101011000000; end
            14'd9097 : begin out <= 64'b0010100101001110001000000100101110011010110101110001111100101100; end
            14'd9098 : begin out <= 64'b1010100000000010101010001011000000010000110011011010100010011000; end
            14'd9099 : begin out <= 64'b0010100011001010001010101111100010101001101000010010001110111111; end
            14'd9100 : begin out <= 64'b0001011000010111100111111100001000100101000111011010001110100000; end
            14'd9101 : begin out <= 64'b0001111001100000001000111111000000101000101101000010000000111001; end
            14'd9102 : begin out <= 64'b0001011100010001001010011111000000100101101011100001110010011011; end
            14'd9103 : begin out <= 64'b0010101000110111001001011001100100101010100000011010011100111010; end
            14'd9104 : begin out <= 64'b1000111010010011101010000101010010101010111110001010100011011101; end
            14'd9105 : begin out <= 64'b1010101001100000101001101010100110101000110101011010011100110101; end
            14'd9106 : begin out <= 64'b1010101110101111000110001111110110101000000100001010000010101101; end
            14'd9107 : begin out <= 64'b0010101010101101000000011110001110101011101010001001111111001001; end
            14'd9108 : begin out <= 64'b0010001110110110001010110100001110101011010101110001111100001110; end
            14'd9109 : begin out <= 64'b1010100101100110001010000011111110100111110010100010101001010000; end
            14'd9110 : begin out <= 64'b1010011111110110100101000111010010101010000010011010001101110001; end
            14'd9111 : begin out <= 64'b1010101101001111101010000010100100101001011011101010011001111100; end
            14'd9112 : begin out <= 64'b1010100110000110001010111011001100101000101011100010011110111100; end
            14'd9113 : begin out <= 64'b1010101000001010101010001010010000101001111100000010001000011111; end
            14'd9114 : begin out <= 64'b1010011111000101001010001110000010101010111010010010011010101110; end
            14'd9115 : begin out <= 64'b1010100110100010101010011110111100100111100000010010101011101010; end
            14'd9116 : begin out <= 64'b0010101110101111101001110101101100101010000110110001111000110101; end
            14'd9117 : begin out <= 64'b0010101101011000001010100110110000100101000000001010101111000110; end
            14'd9118 : begin out <= 64'b0010101001111100101000000101101110101000011001001010101110011100; end
            14'd9119 : begin out <= 64'b1010010110111011100111000010000100101011111100110010100101111100; end
            14'd9120 : begin out <= 64'b0010000101110001001010100001100100100111000010101010100000000110; end
            14'd9121 : begin out <= 64'b0010010110011000001010000111100100101011001111000010101000011110; end
            14'd9122 : begin out <= 64'b1010000011000010101001001010000000101011100100010010100110000011; end
            14'd9123 : begin out <= 64'b0010101111101001000111111001101010101001101111101010100000001111; end
            14'd9124 : begin out <= 64'b0010101000011000001010101010111000100111001111011010011010010101; end
            14'd9125 : begin out <= 64'b1001111100000111001010011110101000011010110110010010101101111010; end
            14'd9126 : begin out <= 64'b1010101000110100101010110011100110101010101100111010000101001110; end
            14'd9127 : begin out <= 64'b0010010001010111101010111101101010011011001011100010000100111010; end
            14'd9128 : begin out <= 64'b1010101101010001001000001000001110100000011010111010011110010011; end
            14'd9129 : begin out <= 64'b0010011111111100001000011101111100101010100100010010000110010000; end
            14'd9130 : begin out <= 64'b1010101010100111000111001100100010101011101001100010010011110101; end
            14'd9131 : begin out <= 64'b0010010000001001001000101010010010011100011100000010101010011101; end
            14'd9132 : begin out <= 64'b0010100010010011000110101010010100100000111001111010100100011111; end
            14'd9133 : begin out <= 64'b1001000001001110101010011000011010011111111111011010100100100110; end
            14'd9134 : begin out <= 64'b1010011110110100001010010111000010100010011001000010010111100000; end
            14'd9135 : begin out <= 64'b0001110001001110001010011001111110101010111000111010101000011011; end
            14'd9136 : begin out <= 64'b0010100100111011001010101110011000100000111011010010000010001100; end
            14'd9137 : begin out <= 64'b0010101101011111101010110001111010011101101001101010100100100110; end
            14'd9138 : begin out <= 64'b1010100000001011001001001110101000101001010111010010100101100000; end
            14'd9139 : begin out <= 64'b0010000010101001001010101010101000100101100111000010101100101010; end
            14'd9140 : begin out <= 64'b0010010110011110101000111100100010100101100100001010100011000100; end
            14'd9141 : begin out <= 64'b0010101000111011001000000001000100100110101000111010011001011110; end
            14'd9142 : begin out <= 64'b1010100111001010001010110101100100101001001000001010101001110011; end
            14'd9143 : begin out <= 64'b1010100100100101001001000000111110101011000110010010101100110101; end
            14'd9144 : begin out <= 64'b1010011010101111101001110000000110101001001000001010100011101001; end
            14'd9145 : begin out <= 64'b1010100000001110001000110011011100100101000010111010100101010101; end
            14'd9146 : begin out <= 64'b0010001001011011001010001011100010010101110010010010011100110111; end
            14'd9147 : begin out <= 64'b0010010100110000101010001101100010101011011010010010010100100011; end
            14'd9148 : begin out <= 64'b1010100110100111001010101101001000101001110011000001100000000010; end
            14'd9149 : begin out <= 64'b0010101101010101001010101011100110101010001000100010101011010100; end
            14'd9150 : begin out <= 64'b1010011110111100000110001001101000100001010000111010100011110111; end
            14'd9151 : begin out <= 64'b1010010101111000001010001010101010100010010010101010100101011111; end
            14'd9152 : begin out <= 64'b0001100100011100001000100000101000101000001110110001110000011000; end
            14'd9153 : begin out <= 64'b1001111001100101000111100001010010100111100011000010100101001001; end
            14'd9154 : begin out <= 64'b1010011010100100101010011110101010101010000111111010001111110101; end
            14'd9155 : begin out <= 64'b1010101101110001001001110111000100101000011010010010100000110110; end
            14'd9156 : begin out <= 64'b0010001000101000101010110001101000101010011111111010011110110101; end
            14'd9157 : begin out <= 64'b0010010001111010101001010001101000101010100110100010011111011000; end
            14'd9158 : begin out <= 64'b0010101011111010001010110100111110101001001001111001100011101111; end
            14'd9159 : begin out <= 64'b0010101001011101101000101101011110100011011010110010101111101101; end
            14'd9160 : begin out <= 64'b1001111011110110001010010101010000011101010001111010101001100101; end
            14'd9161 : begin out <= 64'b0010101010011111001010111011100110101000111101011010010010110101; end
            14'd9162 : begin out <= 64'b1010101101100101100101011010101000100101100000111010101111111001; end
            14'd9163 : begin out <= 64'b1010100000011100101010110110000010101001100000011010011011010101; end
            14'd9164 : begin out <= 64'b1010101111000010100111110100101000101011000110000010101000000011; end
            14'd9165 : begin out <= 64'b1001110011100010101010010100101110011111111101100010010110010110; end
            14'd9166 : begin out <= 64'b0010101001000011001001001111100100100110111100011010100111110011; end
            14'd9167 : begin out <= 64'b0010100101100001001010111111010000101100001111111010100110001110; end
            14'd9168 : begin out <= 64'b1010100011010101101010111001111010101010101000100010101111000111; end
            14'd9169 : begin out <= 64'b0010011011110000101000100011010100101011000010100010100010010000; end
            14'd9170 : begin out <= 64'b0010101000000000100101111000111100101010011100110010001101000100; end
            14'd9171 : begin out <= 64'b1010100010111011001010011100100100100111101000100010100001011001; end
            14'd9172 : begin out <= 64'b0010100010011111001000001000001110100101001001101010101001000111; end
            14'd9173 : begin out <= 64'b0010101000000110001010000011110000100111000001110010101010000111; end
            14'd9174 : begin out <= 64'b0001110100100100001000000111000110100000010101000001110110011010; end
            14'd9175 : begin out <= 64'b0010101101101111100000011110110000011111101111101010101100001100; end
            14'd9176 : begin out <= 64'b0010011010110011101010110001010110100110001010110010100100000100; end
            14'd9177 : begin out <= 64'b1010010011110011001010100011000000100101100001100010000111010011; end
            14'd9178 : begin out <= 64'b0010101110010011101010111111100010101010111000010010100011000101; end
            14'd9179 : begin out <= 64'b1010011011110010101010001010101110100001111110001010101101111001; end
            14'd9180 : begin out <= 64'b0010100101101100001010111110000100100100101100100010101000100100; end
            14'd9181 : begin out <= 64'b0010000010011000101001101111110010101001010001011010100101100011; end
            14'd9182 : begin out <= 64'b0010101010001010001010001111110110100100101111000010011110110010; end
            14'd9183 : begin out <= 64'b1010000101010101101010101110110110011110010100000010011001000110; end
            14'd9184 : begin out <= 64'b1010100000101001001001111000110000101011000010000010100111001011; end
            14'd9185 : begin out <= 64'b1010001100011110001010111011110010101001110110110010100001100011; end
            14'd9186 : begin out <= 64'b1010011101001001101010001100100100011111110001001001010001010010; end
            14'd9187 : begin out <= 64'b0010101101100100101001100100111010101000111000111010101010011000; end
            14'd9188 : begin out <= 64'b1010010111100011001010101001010100100101000111111001001010011101; end
            14'd9189 : begin out <= 64'b1010011101110010101010111010111110101011111010000010010010110101; end
            14'd9190 : begin out <= 64'b0010100010100001101001110111100000100011010101110010011001100011; end
            14'd9191 : begin out <= 64'b0010100110011110001011000011010000101010101011011010100100011111; end
            14'd9192 : begin out <= 64'b0010101111000111101000010010110010101001111000110010001011101011; end
            14'd9193 : begin out <= 64'b1010101001010011001010110111011110100011100101101010010011010000; end
            14'd9194 : begin out <= 64'b0010001110110011101001100101100100100101110100010001111011011100; end
            14'd9195 : begin out <= 64'b1001111101111001001010100010100010100001110100111010100100010101; end
            14'd9196 : begin out <= 64'b0010101000011111001010101111010110101010000100001010001111111000; end
            14'd9197 : begin out <= 64'b0010011000111111101010000100010000011100001100110010000111110010; end
            14'd9198 : begin out <= 64'b0010011001100101101001010110011010101001011010101010010101100010; end
            14'd9199 : begin out <= 64'b1010011110100010101000110011001110101010100111000010101000001101; end
            14'd9200 : begin out <= 64'b0010100010000111101010001101000010011001011101000010100000000010; end
            14'd9201 : begin out <= 64'b0010010001001010001010010111010100101010010100100001110101111100; end
            14'd9202 : begin out <= 64'b0010001000110111101001110001100100101000100000010010101010001100; end
            14'd9203 : begin out <= 64'b1001100100001010000111110111010110101010101101110010100111111011; end
            14'd9204 : begin out <= 64'b1010010111100110100111101001111100011100010001100010101111000000; end
            14'd9205 : begin out <= 64'b0010000011111011101001000100111100100110011101000010101011110000; end
            14'd9206 : begin out <= 64'b0010100000011001101011000010011000100111001101101010100001110110; end
            14'd9207 : begin out <= 64'b1001011001101110101010001111111010101000000010110010011000000011; end
            14'd9208 : begin out <= 64'b0010101101000101101000111001101000101001111100000010101001001011; end
            14'd9209 : begin out <= 64'b0010100110011000101010001100001110101011111100100010001100111011; end
            14'd9210 : begin out <= 64'b1010100101011100001001111011110110101010010100111010001010010011; end
            14'd9211 : begin out <= 64'b1010011001111000101000101010110000100011000100010010100101110010; end
            14'd9212 : begin out <= 64'b1010011111011111001010000011010010101001001011101010100001110111; end
            14'd9213 : begin out <= 64'b0010010010110101100111001101000010101000110000101010100010100111; end
            14'd9214 : begin out <= 64'b0001101001110111101001110100101100100110001110010010100001011001; end
            14'd9215 : begin out <= 64'b0001111000011101001001010101010000101001100010101010100110101011; end
            14'd9216 : begin out <= 64'b1001010100000000101010011110100000101010011100111010100001011111; end
            14'd9217 : begin out <= 64'b1010101000001111001000111011001110100000001001000010101011110100; end
            14'd9218 : begin out <= 64'b0010010100110101101001011010111000100000011111010010001110000010; end
            14'd9219 : begin out <= 64'b0010011110001000001000111110101000100110100000111001110100111000; end
            14'd9220 : begin out <= 64'b1010101110011010101001000001011000100101101101111010011100011111; end
            14'd9221 : begin out <= 64'b0010011110101001100110000100001100101001101011100010101010111001; end
            14'd9222 : begin out <= 64'b0010101011000100001000111000101110101011110111000010001100110110; end
            14'd9223 : begin out <= 64'b1001111000100101101001001110111110100100000110100010000101010100; end
            14'd9224 : begin out <= 64'b1010010010100100001001100110111010101011000110011010101100001110; end
            14'd9225 : begin out <= 64'b1010001001100110101001001000110000100110111101110010110000100010; end
            14'd9226 : begin out <= 64'b0001001100100111101000011000110010101011010111010010100001101111; end
            14'd9227 : begin out <= 64'b1010100110100110000111000110011110100111001111100010000000101111; end
            14'd9228 : begin out <= 64'b1010011100000000101000101101001000101001000000100010011011011011; end
            14'd9229 : begin out <= 64'b1010101101000001101000110111110010100100011001000001110010111111; end
            14'd9230 : begin out <= 64'b0010001011100001100110110110000000100111001001100010101111110000; end
            14'd9231 : begin out <= 64'b1001011101001001101010111000110010100100000011111010100101100110; end
            14'd9232 : begin out <= 64'b0010011111010110101010000000100110101000110110111010010010001001; end
            14'd9233 : begin out <= 64'b0010011011100100001010011011110000011100011111101010100101010101; end
            14'd9234 : begin out <= 64'b0010010010100000101010000000000100101010010001110010011001001001; end
            14'd9235 : begin out <= 64'b1010101010110111101001110011000110101000101010111010100101000101; end
            14'd9236 : begin out <= 64'b1010011111001100001000000010010010101010100101110001111100110010; end
            14'd9237 : begin out <= 64'b1010100001101000101000100110110010101000000101101010100000110101; end
            14'd9238 : begin out <= 64'b1010101001101110101010111011011010011111010101010001110111000000; end
            14'd9239 : begin out <= 64'b1010011111000100001010110110000100100101010100100010101011101101; end
            14'd9240 : begin out <= 64'b0010001000111100001010110010001110100100000011101010010110010011; end
            14'd9241 : begin out <= 64'b1001110011111110000111010101010110101001101001111010100100100000; end
            14'd9242 : begin out <= 64'b1010101001101000001001001100101100101011010011000010001000110110; end
            14'd9243 : begin out <= 64'b1010101100111110000111101101100100100111010010110010000000101100; end
            14'd9244 : begin out <= 64'b0001101101011111001000011101000110101010110111011010010111111100; end
            14'd9245 : begin out <= 64'b0001101101101110001001111011101100100011101101001010101111011110; end
            14'd9246 : begin out <= 64'b1010101010110111001000100010110100100101001001000010101101111110; end
            14'd9247 : begin out <= 64'b1010100001010111001010001110111110101011101100110010100100111110; end
            14'd9248 : begin out <= 64'b1010100111110110000111101101110010100101000001111010101111100101; end
            14'd9249 : begin out <= 64'b1010010101110110101010011000010100101001010010011010100001001100; end
            14'd9250 : begin out <= 64'b0010101100010011001010010110101100101001101101111010101011000010; end
            14'd9251 : begin out <= 64'b0010101101110111001011000010100010100101111000000010011100110111; end
            14'd9252 : begin out <= 64'b0010010001011011101010011011011100011000001000010010100110100000; end
            14'd9253 : begin out <= 64'b0010100010111100101000101011001100100000010001111010011000010100; end
            14'd9254 : begin out <= 64'b1010100000100011100111010111001000101010001010101010000110001000; end
            14'd9255 : begin out <= 64'b1010101010011011001010100101100100010010001000000010011011110101; end
            14'd9256 : begin out <= 64'b1010101010111001001001111100001000100010000111100010011000101111; end
            14'd9257 : begin out <= 64'b1010011001010011001010001000010000011111000101001010001010001100; end
            14'd9258 : begin out <= 64'b0010100110110110101000000100110000101011001001001010101000101111; end
            14'd9259 : begin out <= 64'b1010101111111100101010001010000100011010010110111010101011110001; end
            14'd9260 : begin out <= 64'b0010011010010010000111011111011000011111101100000010100011010001; end
            14'd9261 : begin out <= 64'b0010010100010010101010111101000110100101011101011010011000111010; end
            14'd9262 : begin out <= 64'b0010100100001111101001110011110000101011100011000010001110101011; end
            14'd9263 : begin out <= 64'b0010101001001101001011000011111000101010011000111010100010011010; end
            14'd9264 : begin out <= 64'b1010100010011101101010010100110000101010010100010010101110010110; end
            14'd9265 : begin out <= 64'b1010011011011101001000100110110110101011011101000010100101100110; end
            14'd9266 : begin out <= 64'b1010011111100000101000100101101000100111011100101010100010010101; end
            14'd9267 : begin out <= 64'b0010101010011110101010111001011010100111011111010010000001111101; end
            14'd9268 : begin out <= 64'b0001111111000000001000010100100110100000110101000010101100101011; end
            14'd9269 : begin out <= 64'b1010101001000111001000100111111110101010001000010010010101110001; end
            14'd9270 : begin out <= 64'b0010011101011011101001011110100000100111100110001010100111101101; end
            14'd9271 : begin out <= 64'b1010100110100101001010001001110000100010110011011010000100011101; end
            14'd9272 : begin out <= 64'b0010100100010111001010110100011010100110001011010010011111001001; end
            14'd9273 : begin out <= 64'b1001010111011000001010000110101010101011010100101010101010010011; end
            14'd9274 : begin out <= 64'b0001100100001011000111010000111010101001111101110010101000000010; end
            14'd9275 : begin out <= 64'b1010101010011111001010010011011100100001100110110010000011101100; end
            14'd9276 : begin out <= 64'b0010101101010001101001010011111010101010100000111010100100111000; end
            14'd9277 : begin out <= 64'b1010011101001010001000011011100010100000111001110010010000001101; end
            14'd9278 : begin out <= 64'b0010101110100010101010001011000010100010000010111010100111110010; end
            14'd9279 : begin out <= 64'b1010000011100110100101110100101000101010001111001010101000101001; end
            14'd9280 : begin out <= 64'b1010101011100101001000000100000010100101000011000010101111001000; end
            14'd9281 : begin out <= 64'b1010011001100011101001101101001110100111010011000010011111010110; end
            14'd9282 : begin out <= 64'b1010100100010000001010010011011100100110001011010010100110011111; end
            14'd9283 : begin out <= 64'b1010100011101110001010100010010000101011010110010010011110100101; end
            14'd9284 : begin out <= 64'b1010100011011111101010100110111110011101110000101001010001100100; end
            14'd9285 : begin out <= 64'b1010001010000001001001110110010010100111110111100010100011101010; end
            14'd9286 : begin out <= 64'b1010100100001110001001001010011000101000111110010010100000001111; end
            14'd9287 : begin out <= 64'b1010101000010100101001001011010000100111010111111010100111110110; end
            14'd9288 : begin out <= 64'b1001011101110100001010110010001000101001101011110010100001011010; end
            14'd9289 : begin out <= 64'b0010011111101111100110011011001100001101100010010010010011010001; end
            14'd9290 : begin out <= 64'b0010101001111111101010100100011000100111100010100010100110110000; end
            14'd9291 : begin out <= 64'b1010011101000010101010000000100110101001001110101010011100010111; end
            14'd9292 : begin out <= 64'b1001010110111100001010101000001110101000100000000010100101010101; end
            14'd9293 : begin out <= 64'b1010100001000111100111000100101110011001110010010010101110010100; end
            14'd9294 : begin out <= 64'b0010001011000110101000001110010000101011011111110010100011110101; end
            14'd9295 : begin out <= 64'b0010011100010000101010010110101100100110010100000010101110110010; end
            14'd9296 : begin out <= 64'b0010100011110001000110100010000110101010101000111010100011111010; end
            14'd9297 : begin out <= 64'b1010011001000110101010101100010110011111011000111010010111010011; end
            14'd9298 : begin out <= 64'b0010100101011011001010110101010000101000111101010001011010110001; end
            14'd9299 : begin out <= 64'b1010010000111101100101011000001000100100110011111010101110100110; end
            14'd9300 : begin out <= 64'b0010100101001010101010100001101110011101010100011010000000111001; end
            14'd9301 : begin out <= 64'b0010010110101100001000110100000110100101011100000010001010010000; end
            14'd9302 : begin out <= 64'b0010110001100011001000101101011000011000100011001010010111011010; end
            14'd9303 : begin out <= 64'b1010011100010011001000101100011100101011000111111010100101001110; end
            14'd9304 : begin out <= 64'b1010011010011100001010101010101110010111110100001010010100001000; end
            14'd9305 : begin out <= 64'b1010100110101000001010110101011110101011010010100010011100001001; end
            14'd9306 : begin out <= 64'b1010011100101100101010001101001000101011010110110010011000000001; end
            14'd9307 : begin out <= 64'b1010100101110011101010001010111100100110000100110010001100011100; end
            14'd9308 : begin out <= 64'b0010101010011001101010001110000100011111010001100010011011001011; end
            14'd9309 : begin out <= 64'b1010000011101001101010111000011010101001110101000010100001111101; end
            14'd9310 : begin out <= 64'b1010001110101101101001110110011110011011111000010010100010010111; end
            14'd9311 : begin out <= 64'b0010000011101011101010011011011110011111100101110010000001001100; end
            14'd9312 : begin out <= 64'b0010100001010000001000101010101110101000101100010010011001000110; end
            14'd9313 : begin out <= 64'b1010101011101100001010000110000000101011010011001010011001011000; end
            14'd9314 : begin out <= 64'b1001101001011100101010000001101100010011111110101010101111010011; end
            14'd9315 : begin out <= 64'b1010100010100101001001111111110100100111011111010010101100001010; end
            14'd9316 : begin out <= 64'b0001100001100101001010111011001110101000000100111010011110011100; end
            14'd9317 : begin out <= 64'b1001100010000111001000011001000010101000110000111010100011001101; end
            14'd9318 : begin out <= 64'b0001100010011010001000101101000100101011000010111001111000111000; end
            14'd9319 : begin out <= 64'b0010100101110110101000110111100000100111100000001010101001010100; end
            14'd9320 : begin out <= 64'b1010100101110000001000001000101100101011001000110010010000011011; end
            14'd9321 : begin out <= 64'b0010101011101001001010001001001100100001010001001010011101101011; end
            14'd9322 : begin out <= 64'b1010001101000010001010010010101110100010011111000010011111101011; end
            14'd9323 : begin out <= 64'b1010100011110111101010101011001000101011010100010010010001011001; end
            14'd9324 : begin out <= 64'b0010100010101111101001010001001000100110110011110010100000100010; end
            14'd9325 : begin out <= 64'b0010011110100011101001110100100000101011100101101010010001110000; end
            14'd9326 : begin out <= 64'b0010100000000111001000110101001110100001100110011001100100110111; end
            14'd9327 : begin out <= 64'b1001011010010111001010110110011100100110001000110010001010010010; end
            14'd9328 : begin out <= 64'b0010010100101100101010010000101100011100100111000010100101110100; end
            14'd9329 : begin out <= 64'b0010100001110001001000001001101100101011100011101010100010011111; end
            14'd9330 : begin out <= 64'b1001010010111100101001001110011010100101001111100010101011101000; end
            14'd9331 : begin out <= 64'b1010001110010111000111011001101010011001001001101010011100010000; end
            14'd9332 : begin out <= 64'b1010100101001100101010001111100000101000110101000010101010010111; end
            14'd9333 : begin out <= 64'b0010011110011111101010100011100010100000110110110001101000100000; end
            14'd9334 : begin out <= 64'b1010100010111010101010100110100100101011100100101010100101111100; end
            14'd9335 : begin out <= 64'b1010101010100111001001111101011000101000000110000010010011100111; end
            14'd9336 : begin out <= 64'b0010100001001101101010110000011000100110100010101010101000011111; end
            14'd9337 : begin out <= 64'b1010001100001010001010011001000000101010110110101010001110011111; end
            14'd9338 : begin out <= 64'b1010010000110111001010001101101100100111010001000010100010111100; end
            14'd9339 : begin out <= 64'b0010011001111000001010100101011110100000011001100010011000000110; end
            14'd9340 : begin out <= 64'b0010101010001011101001111011011110010010001010111010011011000101; end
            14'd9341 : begin out <= 64'b1010101100110001000110111100001010100000111001110001011001111101; end
            14'd9342 : begin out <= 64'b0001110111001100000110001101010000101001011110100010100110111010; end
            14'd9343 : begin out <= 64'b1010000111100000000101011001110110011100010001101001111110101111; end
            14'd9344 : begin out <= 64'b0010000011010010001001101010011100101011110001101010010010101101; end
            14'd9345 : begin out <= 64'b1010011110111111101001111110110110100111100010110010110000001101; end
            14'd9346 : begin out <= 64'b1010100110011011001001011010010110101000010101111001001111001010; end
            14'd9347 : begin out <= 64'b1010100011110101001010010000000000101100010000000010110000011001; end
            14'd9348 : begin out <= 64'b0001000101010001101000110101010110101001111001000010100100011101; end
            14'd9349 : begin out <= 64'b1010101110011010101001000000111000100001010110000010100101011111; end
            14'd9350 : begin out <= 64'b0010100001010100101010011001111100100111011100010010010001010011; end
            14'd9351 : begin out <= 64'b1010100101100101101010101000110100100110100011110010010110111010; end
            14'd9352 : begin out <= 64'b1010100111110110001010101011011010100000100001000010011000000110; end
            14'd9353 : begin out <= 64'b1010100111101011101001111100010010100010010000110010101010001011; end
            14'd9354 : begin out <= 64'b0010000100100000100111000101001000101010110110111001010000100001; end
            14'd9355 : begin out <= 64'b1010100110110111101001001010001000101010000101000010000110011011; end
            14'd9356 : begin out <= 64'b1010100010000101001001110100001010100111100010100010101010101010; end
            14'd9357 : begin out <= 64'b1010101000001011101010101110000100011101111110000010101011110100; end
            14'd9358 : begin out <= 64'b1010100001101110101001101111001010100111100110011001111010001000; end
            14'd9359 : begin out <= 64'b0010101110000010001010000010111000100111100111010010101010001100; end
            14'd9360 : begin out <= 64'b0010100100011011101001101001001110100100110100001010011010100111; end
            14'd9361 : begin out <= 64'b0010100101000010001001011110010110101011110011100010100000110001; end
            14'd9362 : begin out <= 64'b1000110100110100101000110000011010101011111101001010101000111001; end
            14'd9363 : begin out <= 64'b1010010101000011101010000111011110100101110001010010101100011011; end
            14'd9364 : begin out <= 64'b0010100100010001001010110100100000100111011011100010011110101010; end
            14'd9365 : begin out <= 64'b0010100001110011101010011111000000101010011111000010101011001110; end
            14'd9366 : begin out <= 64'b0001100010010010001010011111101010011100000111111010110000010001; end
            14'd9367 : begin out <= 64'b1010010111100010101010110111110000101000111001101010101101111111; end
            14'd9368 : begin out <= 64'b1001110111111110001010100110010100101000010001000010101010100111; end
            14'd9369 : begin out <= 64'b0010101010111101001010111100001010100010000011101001111111101000; end
            14'd9370 : begin out <= 64'b1010101011011110100111010001101110101010101011101010001000110110; end
            14'd9371 : begin out <= 64'b1010101011001011001010011100110100101001111010000010010111100000; end
            14'd9372 : begin out <= 64'b1010100011010110101001110111100110011110001101001010101001000001; end
            14'd9373 : begin out <= 64'b1010011011001001101001101110000010101010000011001010100100110000; end
            14'd9374 : begin out <= 64'b0010100001001010001010100000011100100110010110000010110001000010; end
            14'd9375 : begin out <= 64'b0001111101101011101010010011100110100000000000110010100010100011; end
            14'd9376 : begin out <= 64'b1010101100001110000111001001110100101001011101111001011001110001; end
            14'd9377 : begin out <= 64'b0010011111111101001010111111000000011011110110111010100101010111; end
            14'd9378 : begin out <= 64'b1001111010111001001010010100110100100100001110111010000000011001; end
            14'd9379 : begin out <= 64'b1010001001111111001000100101100100100001100111100010100000011001; end
            14'd9380 : begin out <= 64'b0010001010010111001001101111111110101011111101001001110100100011; end
            14'd9381 : begin out <= 64'b1010101101011100101000001010001110101011100101000010011101011110; end
            14'd9382 : begin out <= 64'b1010101001010000101010110101000100011010000101111010101000000001; end
            14'd9383 : begin out <= 64'b1010011001110000001001110111011010100010101010110010101001100011; end
            14'd9384 : begin out <= 64'b0010100111000000000110001000110110100100000101101010100000101000; end
            14'd9385 : begin out <= 64'b1010011010111100001010010110100000101010001111111010100111111101; end
            14'd9386 : begin out <= 64'b1001111110101111001000101010111000011011110011010010100110110111; end
            14'd9387 : begin out <= 64'b1001101010100010101010110111000000101000010011011010100100001110; end
            14'd9388 : begin out <= 64'b1010000100100111001010011011000000101011100101111010100100001010; end
            14'd9389 : begin out <= 64'b0010101101101100001000010111000010100011010011110001111100100010; end
            14'd9390 : begin out <= 64'b0010101000111010101010101000001000011111110111111001000000000100; end
            14'd9391 : begin out <= 64'b0010010111000100001001000101110010011100101110100010100111111011; end
            14'd9392 : begin out <= 64'b0010101010000001001001110110011000100101111111001010101000101110; end
            14'd9393 : begin out <= 64'b1010100101000011001010001100011110101011011000111010001010000010; end
            14'd9394 : begin out <= 64'b0010100000011110101010001011110100100110100010101010000100001111; end
            14'd9395 : begin out <= 64'b1010010100101001001010010100000100101010000011100010010111101011; end
            14'd9396 : begin out <= 64'b1010000110101001101010100111100010100100100000101010100011011001; end
            14'd9397 : begin out <= 64'b1010100001110111001000101000110000101000101100011001111000000110; end
            14'd9398 : begin out <= 64'b0010010110011001001000010001010110101000010010001010001111000111; end
            14'd9399 : begin out <= 64'b1010101001100100001011000010111100100110010110010010100110010100; end
            14'd9400 : begin out <= 64'b0010010100010001001001100110001100100110101000010001110111101111; end
            14'd9401 : begin out <= 64'b1010011000111110100111111100101100101010111001000001000111100110; end
            14'd9402 : begin out <= 64'b0010100011101011100110101110000010101000110111110010100111110110; end
            14'd9403 : begin out <= 64'b0010100111100000001011000101000110100111011010001010010100001111; end
            14'd9404 : begin out <= 64'b1010010111110000101000010110100100101011000000100001001000010100; end
            14'd9405 : begin out <= 64'b0010011001101000101010111111101000101001001001110010101100101100; end
            14'd9406 : begin out <= 64'b1010010010100110101010110110110110100011111110111010011000001110; end
            14'd9407 : begin out <= 64'b1010101110011000101000001110001100011100011000100010010011001101; end
            14'd9408 : begin out <= 64'b1010100000100001100110000001100000101011011111110010010110111111; end
            14'd9409 : begin out <= 64'b0010011001101001001010011110000110100101111101010010100101100100; end
            14'd9410 : begin out <= 64'b0010000100010001001001100100101000100000100010110010101001000010; end
            14'd9411 : begin out <= 64'b0010101010110000001010010011111010100101110010100010100000100000; end
            14'd9412 : begin out <= 64'b1010101001111101101001111111000110101011010110111010011110100010; end
            14'd9413 : begin out <= 64'b0010100000001111100110110110010110101100000101010010000011001110; end
            14'd9414 : begin out <= 64'b0010100111101001101010101110100110101100001001011001010110100111; end
            14'd9415 : begin out <= 64'b1010100100101110101000110111010000011010110101101010100000010101; end
            14'd9416 : begin out <= 64'b1010100010100010101001110001000110101001001000110010010110010101; end
            14'd9417 : begin out <= 64'b1010101110010010001010110011100110101000010011100010101110101101; end
            14'd9418 : begin out <= 64'b0010100110100101101001111110111100100110000010011010101001101100; end
            14'd9419 : begin out <= 64'b0010011111011111001001100000100110101000001110111010011110110110; end
            14'd9420 : begin out <= 64'b0010010101000011101011000001111110100011010101101010011010000010; end
            14'd9421 : begin out <= 64'b1010100111111101001010011001011000101011110110101010101101100100; end
            14'd9422 : begin out <= 64'b1010101011000011101001000110011100101011101111010010101001110011; end
            14'd9423 : begin out <= 64'b1010010111010010101010000010010010001000111000110010110000000011; end
            14'd9424 : begin out <= 64'b0010100011110111001001001001110010100111011100001010101011101001; end
            14'd9425 : begin out <= 64'b1010100011011101101010101110001000101011000101111010000000100010; end
            14'd9426 : begin out <= 64'b0010010011101011001010000100010100101010110001010010010100100101; end
            14'd9427 : begin out <= 64'b0010101101111110001010010101101010101001001111000010100001111100; end
            14'd9428 : begin out <= 64'b0010010000010111101010010011001010100111100100110010100100011001; end
            14'd9429 : begin out <= 64'b1010011001011011001001110111111110100110101110100001111111000100; end
            14'd9430 : begin out <= 64'b0010011010110000001010111100101110101011011100000010100000110001; end
            14'd9431 : begin out <= 64'b1010001011011000101010000111100010101011110011001010010010011101; end
            14'd9432 : begin out <= 64'b1001110111100111001001110000101100101011101010110010101000010100; end
            14'd9433 : begin out <= 64'b0010100111100100001010011110010110100110101011010010100111000110; end
            14'd9434 : begin out <= 64'b1010001011010001001010011011110110101010011010111010100011100011; end
            14'd9435 : begin out <= 64'b1010101111100100001001000011100000100111101110100010100001110010; end
            14'd9436 : begin out <= 64'b1010100000001100001001100000000010100100101100101010101011110101; end
            14'd9437 : begin out <= 64'b1010010011110110101001101111100010101011100111101010011001000001; end
            14'd9438 : begin out <= 64'b1010010000110110101010101111010100101011010111011010100111010011; end
            14'd9439 : begin out <= 64'b0010100011010110001010110010000100100101110100001010101001000111; end
            14'd9440 : begin out <= 64'b0010101011001110101010100111000100100111010001011001110101101010; end
            14'd9441 : begin out <= 64'b1010100111111010001010010111101000011011000100111010000000000110; end
            14'd9442 : begin out <= 64'b0010010100101011101010101010010100101000000001010010101111010101; end
            14'd9443 : begin out <= 64'b1001111010010011100110001010110000101011110010110010000101110110; end
            14'd9444 : begin out <= 64'b1010000010111010000110010101100000011010010100000010100001000111; end
            14'd9445 : begin out <= 64'b0010001000101100001001111111000000101011101101011010100100101101; end
            14'd9446 : begin out <= 64'b0010010010101101101010001000101010101011100100010001001110100110; end
            14'd9447 : begin out <= 64'b0001101000101110001001100110111100011010101110001010101000010100; end
            14'd9448 : begin out <= 64'b1010101100000000101010001000111000101011101001110001111110011100; end
            14'd9449 : begin out <= 64'b0010100100100011001010100001110110011010000010110010000101101101; end
            14'd9450 : begin out <= 64'b0010010111001011001001000001000010101001001001010010010000100010; end
            14'd9451 : begin out <= 64'b0010100100011001101010011010101000100100000000100010100110110110; end
            14'd9452 : begin out <= 64'b0010100100001001101000010101101110101000001010000010001111100001; end
            14'd9453 : begin out <= 64'b0001110111100111001001011000100010100111101100101010100101110101; end
            14'd9454 : begin out <= 64'b1010101110111011101010100010101010101011001001110010100100101011; end
            14'd9455 : begin out <= 64'b0001100111111100001010011101100110100100010000010010001000000101; end
            14'd9456 : begin out <= 64'b1010001110000010100110111100000100100000011000001010100000011111; end
            14'd9457 : begin out <= 64'b1010100101110110001010101100110000100101011001011010000111110111; end
            14'd9458 : begin out <= 64'b1010001000101100001001011111001100001001001111111001110011100101; end
            14'd9459 : begin out <= 64'b0010100011111011101010101010101100100101110100100001111100101111; end
            14'd9460 : begin out <= 64'b0010011011100000001000101001100110101000001001000010100010010111; end
            14'd9461 : begin out <= 64'b0010100101000110001011000001100010100000111110111001011101011011; end
            14'd9462 : begin out <= 64'b0010101011111011001010100001011010101011110011100010101000001100; end
            14'd9463 : begin out <= 64'b1010010111010010101010001110000010101001111100001010100111111001; end
            14'd9464 : begin out <= 64'b1001111101111010101001111101010010101000011111011010101001111010; end
            14'd9465 : begin out <= 64'b0010101100001011001010011011111010101000110101010010101010111010; end
            14'd9466 : begin out <= 64'b1010101010100000001000010111000000101010110111011010101000101101; end
            14'd9467 : begin out <= 64'b0010010101100100101010010011000010101011001110110010100001101010; end
            14'd9468 : begin out <= 64'b1010100100110010001001101010100000100100001110010001101101010010; end
            14'd9469 : begin out <= 64'b1001110000011100101010010111111100100110100111101010001011000111; end
            14'd9470 : begin out <= 64'b0010100001010110000111000101001000100100110000101010011011010100; end
            14'd9471 : begin out <= 64'b0010100101111111101000001010100000100110001010001010011100001001; end
            14'd9472 : begin out <= 64'b1001100110110001101010100001100010101010011110010010100001010110; end
            14'd9473 : begin out <= 64'b1010011011110000101001001101110000100011000110001010100010111111; end
            14'd9474 : begin out <= 64'b1010010110000100001001100001010000100101000111001010010011010001; end
            14'd9475 : begin out <= 64'b0010010100111011101010000001111100100100010110101010010100011010; end
            14'd9476 : begin out <= 64'b0010100000000000101000010111100100101001111011100010000101100010; end
            14'd9477 : begin out <= 64'b1010101001000000001010000001011000100001111000101010100000011011; end
            14'd9478 : begin out <= 64'b0010101000010000001010110001101100101001110010011010011111001110; end
            14'd9479 : begin out <= 64'b1010101101111111101001110010001110101011000101101010101000110010; end
            14'd9480 : begin out <= 64'b1010100010101001001010011000100000101011110101000010001111101010; end
            14'd9481 : begin out <= 64'b0010010110100101101010101011010100100000111001101010010111010100; end
            14'd9482 : begin out <= 64'b1010010010110110001001001001001000011010111111010010100000011111; end
            14'd9483 : begin out <= 64'b1010010111000111001001011111010000010011000000000010101010011101; end
            14'd9484 : begin out <= 64'b0010101011100100001010100001000110100101111110000010000110100000; end
            14'd9485 : begin out <= 64'b1010011011101111101000010101010010100101100001101010010100100000; end
            14'd9486 : begin out <= 64'b1001110111100001001010011111011110100110000110110010101000001111; end
            14'd9487 : begin out <= 64'b1010100101100011101010111100101100101001011010011010101100101001; end
            14'd9488 : begin out <= 64'b0010100010110000101001110001000100100110100001111010100000011100; end
            14'd9489 : begin out <= 64'b0010010011101111001001000100011100101001110111110010101011011101; end
            14'd9490 : begin out <= 64'b1010010000001100000110010001101010101011011100110010101001101111; end
            14'd9491 : begin out <= 64'b1010010010010001101010010010111100101010110011010010001110010101; end
            14'd9492 : begin out <= 64'b0010100110111110101001000110010100101010111000101010101011000101; end
            14'd9493 : begin out <= 64'b1010010100110000101010010111001100100110111010100010000011111001; end
            14'd9494 : begin out <= 64'b1010100010100100001001000100011110101010111100111010101111011111; end
            14'd9495 : begin out <= 64'b0010101000010011101010100000010010100110100011100001111011101000; end
            14'd9496 : begin out <= 64'b1010100101101110001010101000001110100011101010001001111010111001; end
            14'd9497 : begin out <= 64'b0010010110001001001001000100110100101000100101011010100000011100; end
            14'd9498 : begin out <= 64'b1010010100101100101010011000111110011100010001101010101111000101; end
            14'd9499 : begin out <= 64'b1010100101110011101010101000111000011100111100010010100001010110; end
            14'd9500 : begin out <= 64'b1010001101100001001010100001010110100001100101110010010101001000; end
            14'd9501 : begin out <= 64'b1010010101010010101000000011010000101000111001000010010011010101; end
            14'd9502 : begin out <= 64'b1010000011110011101010110111011000100000011000011010100111001101; end
            14'd9503 : begin out <= 64'b1010100011011101101001110111010010100100001000111010100010100011; end
            14'd9504 : begin out <= 64'b0010100101111001001000111001111110011101101000001010101000101001; end
            14'd9505 : begin out <= 64'b0010101010001110001010100101000000101001010111000010001101011011; end
            14'd9506 : begin out <= 64'b1010000001001101001010110000000110101000100101101010100100001001; end
            14'd9507 : begin out <= 64'b1010101000111000001010111101001000100101001100000010101101101100; end
            14'd9508 : begin out <= 64'b1010010111111001001010011010000110100101101001011010010010011100; end
            14'd9509 : begin out <= 64'b1010100011010011101010001111001110101010100100011000110101000110; end
            14'd9510 : begin out <= 64'b0010101100011010100111100101010010011101101110010010100100101110; end
            14'd9511 : begin out <= 64'b1010100101110011001010010111000000101000011001111010010101000011; end
            14'd9512 : begin out <= 64'b1010101001000111000111110001100110101011011010111010010100000010; end
            14'd9513 : begin out <= 64'b0010101010111110001010111100001100101000011101011010100100111010; end
            14'd9514 : begin out <= 64'b0010110000000111001001100110000100100110000101011010101010011100; end
            14'd9515 : begin out <= 64'b1010101010000001001000101011010000100111010010010010011001100011; end
            14'd9516 : begin out <= 64'b0010011011010011101010101100000100101011001101110010011001011101; end
            14'd9517 : begin out <= 64'b1010010011000001101010110010011100100111110110100010011100001010; end
            14'd9518 : begin out <= 64'b1010101001011110101010000111111100101001011010011010101111001110; end
            14'd9519 : begin out <= 64'b0010100000011101001010000001010100100100111100011010100011011011; end
            14'd9520 : begin out <= 64'b0010100110011111001010100100100110101001001111010010100110001101; end
            14'd9521 : begin out <= 64'b1010100111000111101010010111101010100110000000111010101001000000; end
            14'd9522 : begin out <= 64'b0010010011011000001001001110001110101010100011110010010010110101; end
            14'd9523 : begin out <= 64'b1010010010001011101010100101011100100010101101000010100101010110; end
            14'd9524 : begin out <= 64'b0010101010000101101010011011110000011011111001000010101101011110; end
            14'd9525 : begin out <= 64'b0001110011101001000000000010100100101011100101110010000110001010; end
            14'd9526 : begin out <= 64'b0010101101100010001010011111010010011001101001101010011011001111; end
            14'd9527 : begin out <= 64'b1010100110011011001010001001100100101010010110101010001010100111; end
            14'd9528 : begin out <= 64'b0010011000010111101001101101010010100100001010101010100101100000; end
            14'd9529 : begin out <= 64'b0010011100000111101001101010011100101011100101011001110101010010; end
            14'd9530 : begin out <= 64'b0001110001001111101010111001010010100101110001001010100000100111; end
            14'd9531 : begin out <= 64'b0001110101101111101010000101100100101000110010111010000111111011; end
            14'd9532 : begin out <= 64'b0010100001100111100101111111101010100110001010101010100101111101; end
            14'd9533 : begin out <= 64'b0010101001110010000101100111110000101011100111110010101111000000; end
            14'd9534 : begin out <= 64'b1010011001111101101010100110010010100111000010110010010111110010; end
            14'd9535 : begin out <= 64'b1010101101100010100111100100110000100000000100000010101011101101; end
            14'd9536 : begin out <= 64'b1010100010111011101001100110011000100111001001110010100110110100; end
            14'd9537 : begin out <= 64'b0001110000001111101010100011010010100011110001110010101110110011; end
            14'd9538 : begin out <= 64'b0010010110100101101000101111001100100110100001010010001101100101; end
            14'd9539 : begin out <= 64'b1010010000111100001001000011100100101001000011011010101101001111; end
            14'd9540 : begin out <= 64'b0010001101101001001010010010011010101001110011110010100000101011; end
            14'd9541 : begin out <= 64'b0010010111011011101010100111011000100111100100010010000011000111; end
            14'd9542 : begin out <= 64'b1010001111100011001010010011000110100101001000000010000001110000; end
            14'd9543 : begin out <= 64'b0010100111000101101010011010001010101010010000101010101111101011; end
            14'd9544 : begin out <= 64'b0010010110001011001010000001111000101011001001111010011000011011; end
            14'd9545 : begin out <= 64'b0010101100110000001001100000000010101000011001001001100111010110; end
            14'd9546 : begin out <= 64'b0010100000011100001010001000011110100011111001001010011100010101; end
            14'd9547 : begin out <= 64'b0010000001111111001010101001011110100111111000001010100011010000; end
            14'd9548 : begin out <= 64'b0010101000100010001001111000000100101001110000101010001000010101; end
            14'd9549 : begin out <= 64'b0010101011001011101000111011001100100111111111110001110100100101; end
            14'd9550 : begin out <= 64'b0010000010000000101010101010000010010100101000000010000100001110; end
            14'd9551 : begin out <= 64'b1010011111101101001010110000001100101000011010000001111010111011; end
            14'd9552 : begin out <= 64'b0010101000001111101000001110001110101000111001110010011100111011; end
            14'd9553 : begin out <= 64'b0010101101001100000101101111101000100101111011110001000100111000; end
            14'd9554 : begin out <= 64'b0010100011101110001001111000101010101011110100110001111111111000; end
            14'd9555 : begin out <= 64'b1010100110010000101010000011000010011001011110101010100111111011; end
            14'd9556 : begin out <= 64'b1010101110010101001010000011111010100111011111001010100010011100; end
            14'd9557 : begin out <= 64'b1010100001010101101001010010000100101001000000011010011000100001; end
            14'd9558 : begin out <= 64'b0010010101100111001000000010111110101000101110100010101101111000; end
            14'd9559 : begin out <= 64'b0010101101111100101001100111110110101011010011101010100000110110; end
            14'd9560 : begin out <= 64'b1001101010110101000100001001101100011100110011100010010010111001; end
            14'd9561 : begin out <= 64'b1010100010110010001010110110001010101000111101100010000000001010; end
            14'd9562 : begin out <= 64'b0010000011011110101010001000101010101010110100011010001100001001; end
            14'd9563 : begin out <= 64'b1010011010010010001010000100111110100001110001111001100101010110; end
            14'd9564 : begin out <= 64'b0010000111100111001010101100010000101001000010111010100011111110; end
            14'd9565 : begin out <= 64'b1010000000000111101010101110101110101011101011010010101010100010; end
            14'd9566 : begin out <= 64'b1010101000011100001001100110001100100111110010001010101011101110; end
            14'd9567 : begin out <= 64'b1010100111101111000110001000110010100010000001110010101101000100; end
            14'd9568 : begin out <= 64'b1010101111110010001001100000011010101011000100010010101000100111; end
            14'd9569 : begin out <= 64'b0010010100100100101001011001111000101000011010100010011101011010; end
            14'd9570 : begin out <= 64'b1010101001111111101010011010110110101010010001111010101101010111; end
            14'd9571 : begin out <= 64'b1001111011111101001010011111001010100111100010010001110111000001; end
            14'd9572 : begin out <= 64'b0010101011000101000111001010001000101000110110011010100100100010; end
            14'd9573 : begin out <= 64'b1010100101001001100110000111100000100101100111111010101101101101; end
            14'd9574 : begin out <= 64'b0010010101101000100110000010111100101000111011110010100001011100; end
            14'd9575 : begin out <= 64'b0010010001010000001001011010111100100100100010111010011101101010; end
            14'd9576 : begin out <= 64'b1010010110111011001010011111000110101011001100010010100101010011; end
            14'd9577 : begin out <= 64'b1010010110000010101001110100100010101010100101000010000101100000; end
            14'd9578 : begin out <= 64'b0010100100010111101001100110000010101000011110000010100110101110; end
            14'd9579 : begin out <= 64'b0010011010101111001010010000100100101001110010001010100001010011; end
            14'd9580 : begin out <= 64'b1010011010010100101010100011100100101000101101111010100000110000; end
            14'd9581 : begin out <= 64'b0010001000101111001001111010111010101001110111110010000011010101; end
            14'd9582 : begin out <= 64'b0010011000001010101010111101010110101001111010000010000001100101; end
            14'd9583 : begin out <= 64'b1010100100001010101010110110100100100011100110110010010000001100; end
            14'd9584 : begin out <= 64'b0010100100100101101010011001101010100111011100110010010100110011; end
            14'd9585 : begin out <= 64'b1010100001111111100110111010011110100010110111001010010100011001; end
            14'd9586 : begin out <= 64'b0010010100111001101001001100010110100111101100001010010101000011; end
            14'd9587 : begin out <= 64'b0010000011011100101010011111101100100100110001101010011001100011; end
            14'd9588 : begin out <= 64'b0010100001110011101001010010111010101011011010001010101010110101; end
            14'd9589 : begin out <= 64'b1010011101110101001010101100100100101000111100110010011110011011; end
            14'd9590 : begin out <= 64'b0010101000010011101000111001101000101011000111001001111010011101; end
            14'd9591 : begin out <= 64'b1010100100000100000101011111101100101010000110111010100010111010; end
            14'd9592 : begin out <= 64'b1001110110101001101001000110101000100101110100011010011001010111; end
            14'd9593 : begin out <= 64'b1010001101000110001010110100001100101001100000101010011100100111; end
            14'd9594 : begin out <= 64'b0010100101100100101010000010101000101001000111111010001001111100; end
            14'd9595 : begin out <= 64'b1010100011111010101000011010010010100111010010100001110010110001; end
            14'd9596 : begin out <= 64'b0001011101010000001001110100111110100110011011010010101100001011; end
            14'd9597 : begin out <= 64'b1010000111000100001010000000100100101001101010110010100000110101; end
            14'd9598 : begin out <= 64'b1010011110010101101010000010111110011101110101111010101101100111; end
            14'd9599 : begin out <= 64'b1010000000110001001010101011000110100111111010100010100101101000; end
            14'd9600 : begin out <= 64'b0010100011110011001010111001101000101001100101111001111111001010; end
            14'd9601 : begin out <= 64'b1001111110110111000101000001111000100111100111001010101111101011; end
            14'd9602 : begin out <= 64'b1010010001101100001010010110010000100000100100100001100101001000; end
            14'd9603 : begin out <= 64'b1010000100001111001001011001110000101001100010110001111101100111; end
            14'd9604 : begin out <= 64'b1010100010001100001010010110001110100010010101100010011011111111; end
            14'd9605 : begin out <= 64'b0010000100011011100111011010100000101000010101101010101001000000; end
            14'd9606 : begin out <= 64'b1001111110010100001010011001111100100110010100101001101111101000; end
            14'd9607 : begin out <= 64'b1010000010100111001001110110000100101001001101110010100110110000; end
            14'd9608 : begin out <= 64'b1010010001111011101010100101011010101011101010011010100001010101; end
            14'd9609 : begin out <= 64'b0010101001000011101000101110000010101001011100111010100011001100; end
            14'd9610 : begin out <= 64'b1010100111011100101000101111110100101001011111100010100010011111; end
            14'd9611 : begin out <= 64'b1010001100010110100101001101010010101001000011110010011010100101; end
            14'd9612 : begin out <= 64'b0001110110001110001000001100011000100110010010100010010000001010; end
            14'd9613 : begin out <= 64'b1010001010000100001010010101110100100001001111000010011010100011; end
            14'd9614 : begin out <= 64'b0010101100010100100110101110001100100100000010000010010000100101; end
            14'd9615 : begin out <= 64'b0010001111010110001010010010111000101000100111000010010010011011; end
            14'd9616 : begin out <= 64'b0010000010001100000111010011111110011101010100011010011000101110; end
            14'd9617 : begin out <= 64'b1010010101000011101000011111110100011010100000010010110000010001; end
            14'd9618 : begin out <= 64'b0001111010001001001001101111101100011110001100001010100010000011; end
            14'd9619 : begin out <= 64'b0010100101011010001000101100100010101011010001011010010111110001; end
            14'd9620 : begin out <= 64'b0010010101000000001001000110010000101001010100111010001100000110; end
            14'd9621 : begin out <= 64'b0010011101010100101001100110111110101000001011100010011101001101; end
            14'd9622 : begin out <= 64'b0010011100010010001010100000100110101011111100010010100011000011; end
            14'd9623 : begin out <= 64'b1010100001111110001010100100010110100101001000000010010100100101; end
            14'd9624 : begin out <= 64'b1010011011011010101010000110111100101000010101110010100010101000; end
            14'd9625 : begin out <= 64'b0010001000011110101010100001011100100001111001010010001000111000; end
            14'd9626 : begin out <= 64'b0010101000111000000111000111101010100000011000010001101000010111; end
            14'd9627 : begin out <= 64'b0010100000100001101010110100010010101010111110000001111001000110; end
            14'd9628 : begin out <= 64'b1010011111010110101001111110111010100101000000011010011111010001; end
            14'd9629 : begin out <= 64'b1010010111100110001000011100000110101001100000111001110100000011; end
            14'd9630 : begin out <= 64'b0010000101001011001000001010000010100011011101110010101010100000; end
            14'd9631 : begin out <= 64'b0010101011011110101010010000001010011100110000111010011000111110; end
            14'd9632 : begin out <= 64'b0010011110100011101010101010110100100101011011001010011011000010; end
            14'd9633 : begin out <= 64'b0010000000111010101010100101100010101000010111000010001111100001; end
            14'd9634 : begin out <= 64'b0010011011111101100101101011000110101010010100111010010011100000; end
            14'd9635 : begin out <= 64'b0010100111010001101000101111001010101000111111001010101010111001; end
            14'd9636 : begin out <= 64'b0010001100000101001010011110000100100101011010110010100101111000; end
            14'd9637 : begin out <= 64'b0010100010101010101010011100100010100110101110000001110100110011; end
            14'd9638 : begin out <= 64'b1010011010100111101010100110111110100100110011011010100010001100; end
            14'd9639 : begin out <= 64'b1010101110100110001010111011101110101011010000000010011111001010; end
            14'd9640 : begin out <= 64'b1001101100001110001000000100110100011101010100100010100010101011; end
            14'd9641 : begin out <= 64'b0010010001011110101001011011101000101011110000110010001101011010; end
            14'd9642 : begin out <= 64'b1001111110100111101010110001111110101010110101000010101110101010; end
            14'd9643 : begin out <= 64'b1010101111010011101010000011111000100111101101011001100001011100; end
            14'd9644 : begin out <= 64'b1010100110000010100111100000101000101010100111001010101111010000; end
            14'd9645 : begin out <= 64'b1010101110010111000110010110110110101001001101011001011000000110; end
            14'd9646 : begin out <= 64'b0010001000011110001010110001110100101000011101101010100000111101; end
            14'd9647 : begin out <= 64'b1010011001001111001010010100001010101000111011100010011000111100; end
            14'd9648 : begin out <= 64'b1010100010001001001001010100101010101001001100010010000111001000; end
            14'd9649 : begin out <= 64'b0010101010000111101010001111011000101000101101001010010111011011; end
            14'd9650 : begin out <= 64'b0010010011010100101001000010110010101000101110000010001001011101; end
            14'd9651 : begin out <= 64'b1010100010101110101010111100001110101000110010110010101011000010; end
            14'd9652 : begin out <= 64'b1010010110010110101010111010111000101010011010111010100100010100; end
            14'd9653 : begin out <= 64'b1010101000010100001000000000010000101010010010000010100001000100; end
            14'd9654 : begin out <= 64'b1010000110111000001010001100001110100111001100100010100111010000; end
            14'd9655 : begin out <= 64'b1010101110110000001010000101011010100100111100010010011100001001; end
            14'd9656 : begin out <= 64'b0001101001010010101010000011000010100011111111110010101110101111; end
            14'd9657 : begin out <= 64'b1010010110011101001000001010000100101010010101000010011111111010; end
            14'd9658 : begin out <= 64'b1010010011011101001010001111011100101011010110000010001101010100; end
            14'd9659 : begin out <= 64'b0010011000100100001001110011111110011110000100000010010111111001; end
            14'd9660 : begin out <= 64'b1010100011000111001001100010100110011110011110010010101000110011; end
            14'd9661 : begin out <= 64'b0010011101100000001000100011010000010101010000001010100101010000; end
            14'd9662 : begin out <= 64'b0010001101011100001001010011110010101010000010101010101010001011; end
            14'd9663 : begin out <= 64'b0010100011001100001001110100101100100000110110001010101001011111; end
            14'd9664 : begin out <= 64'b0001101100100111001010011111111110101010101110001010011000110001; end
            14'd9665 : begin out <= 64'b0010100000101101101001001011110010101000101110111010101100111010; end
            14'd9666 : begin out <= 64'b1010100111000100001010011100000100101000110000010010000011111000; end
            14'd9667 : begin out <= 64'b0010001101010111001010110001000010100110000110010010100011010101; end
            14'd9668 : begin out <= 64'b0010101000111000101001010010000010101011101111110010011110110101; end
            14'd9669 : begin out <= 64'b1010100010010011001010100011100000011001000010100010100000010001; end
            14'd9670 : begin out <= 64'b1010100100000011001010010011110110101000100011001010001000101011; end
            14'd9671 : begin out <= 64'b1010100011101111101010100011010010011011011011100010101111001101; end
            14'd9672 : begin out <= 64'b1010010011110101001001100110011000101010110000110010011010001111; end
            14'd9673 : begin out <= 64'b0010101110101011101000100010101100101010101101111010010011011101; end
            14'd9674 : begin out <= 64'b1010101011011010101001001001010010101011111000010010100011011010; end
            14'd9675 : begin out <= 64'b1000110010010111001001011011111100100101111001101010010101111000; end
            14'd9676 : begin out <= 64'b1010101101000000001010100001110010101011101110110010000010001110; end
            14'd9677 : begin out <= 64'b1001111100010101001010111010000110100100001011011010100010100111; end
            14'd9678 : begin out <= 64'b1010100100010101001001010111101110101010011110110010010011101010; end
            14'd9679 : begin out <= 64'b0010001010001000101010111000110000100100000011001010011110010001; end
            14'd9680 : begin out <= 64'b1010101110111001100111101100001110101001100000000010100100111001; end
            14'd9681 : begin out <= 64'b1010100011001001101010100101010000101000101000101010100101111000; end
            14'd9682 : begin out <= 64'b1010101001110111101010011010010110101011100111110001100011001010; end
            14'd9683 : begin out <= 64'b1010101111001010001010101001111000100001110000110010010011000101; end
            14'd9684 : begin out <= 64'b1010000001110001101010110011111010101001100111010010100100111100; end
            14'd9685 : begin out <= 64'b0010000010010111001010010010111100101001100111110010101010000111; end
            14'd9686 : begin out <= 64'b0010011001110110101001001100100000100000101000111010010010111101; end
            14'd9687 : begin out <= 64'b1010000010011100101001010001110000101000000001011010100010010100; end
            14'd9688 : begin out <= 64'b1010101010111001101001101000011010100011000010111010100101111011; end
            14'd9689 : begin out <= 64'b0010011011110011001010110100101000101010010011100010100101001010; end
            14'd9690 : begin out <= 64'b1010100101010011001010011001111110101010001010110010011100100001; end
            14'd9691 : begin out <= 64'b1010100110001100001000001010010010101010111010000010101111000100; end
            14'd9692 : begin out <= 64'b1010101010010101000111001001101000100100010111010010011000011111; end
            14'd9693 : begin out <= 64'b1010100001000001001010110100101000100000000001010010001001111011; end
            14'd9694 : begin out <= 64'b1010100011101111001010111100001100100010010100101010011111110010; end
            14'd9695 : begin out <= 64'b1010011111100100101001010101000000101000100001010010101101010110; end
            14'd9696 : begin out <= 64'b1010101100011100101010101101111010011100011011000010010111011001; end
            14'd9697 : begin out <= 64'b0010101000001101001010111010110100100101000000111010011000100101; end
            14'd9698 : begin out <= 64'b1010100010011010000111011011000100101010111100011010010011011111; end
            14'd9699 : begin out <= 64'b1010100100101011001001111101100100100110001111101000101110111110; end
            14'd9700 : begin out <= 64'b0010101101100111101010101011011000101000000111011010101010101000; end
            14'd9701 : begin out <= 64'b1010010111010010001001111101111110100100010100001010000001101100; end
            14'd9702 : begin out <= 64'b1010101001100101001000010000111110101011010011100010100011111111; end
            14'd9703 : begin out <= 64'b0010100101011011101010011011001000100110001101001010101001111101; end
            14'd9704 : begin out <= 64'b0010011101101010001000000111000010100011111001000010010111001001; end
            14'd9705 : begin out <= 64'b1010011011011111101001100110100000101011111100111010100101100101; end
            14'd9706 : begin out <= 64'b0010101010100101001010011001110010100000100011111010101100111100; end
            14'd9707 : begin out <= 64'b1010100101001100001010010011101100101011010111001010001000000110; end
            14'd9708 : begin out <= 64'b1010100011001100100100111111101110101001001100001010001110000111; end
            14'd9709 : begin out <= 64'b0010100000011111001000001101001100101000011110001010101100011111; end
            14'd9710 : begin out <= 64'b1010001111101101001010011011011110101011001000111010101110100110; end
            14'd9711 : begin out <= 64'b0010000001001100001010001001010000101011110110010010011111101000; end
            14'd9712 : begin out <= 64'b1010101010011110100111100011010110010100011101010001101001100000; end
            14'd9713 : begin out <= 64'b0001011111011001001001100010100100101000110101011010011110010010; end
            14'd9714 : begin out <= 64'b1010101111001000101010001010100000011100010110101001111100100110; end
            14'd9715 : begin out <= 64'b0010101001101100001001101110011110011001000001100010101010011110; end
            14'd9716 : begin out <= 64'b0001110101000000001001010100000000100101101101000010100001111011; end
            14'd9717 : begin out <= 64'b0010100101010101101001000101100010101011000000110010101110101110; end
            14'd9718 : begin out <= 64'b1010101100001100001001101010001110100111001101011010101101100000; end
            14'd9719 : begin out <= 64'b0010011010011010101001011000100010100110010111000010101101111111; end
            14'd9720 : begin out <= 64'b0010100100000001001010111010111100100001100011100010000011000011; end
            14'd9721 : begin out <= 64'b1010000000011100101000001110010110100001101001111010101111111011; end
            14'd9722 : begin out <= 64'b0010101111101001101001011000000000101011010101100010011011110101; end
            14'd9723 : begin out <= 64'b0010101100001010001010110010111100011110101110001010100111110001; end
            14'd9724 : begin out <= 64'b1010011010000000101010100111101110101001100100010010010101100001; end
            14'd9725 : begin out <= 64'b0010101010000001100110101100111110101010000110100001100111000100; end
            14'd9726 : begin out <= 64'b0010100110010001101010011011110000101011001001100010001010111111; end
            14'd9727 : begin out <= 64'b0001110011100011001010010110000000101100001001001010100111000011; end
            14'd9728 : begin out <= 64'b0001000000111001101001110110010100101011111111001010001100010100; end
            14'd9729 : begin out <= 64'b0010000111010000001001110111100000101000000111010010011110011010; end
            14'd9730 : begin out <= 64'b1001111010101010001010001011110110101001111100011010101100001100; end
            14'd9731 : begin out <= 64'b0001101011001010101001100001011100100001110001010001110111000101; end
            14'd9732 : begin out <= 64'b0010101001001010101001100001111000011101100001000010010101010010; end
            14'd9733 : begin out <= 64'b0010011010101101001001011011100110100000111101110001001011111000; end
            14'd9734 : begin out <= 64'b0010100000111001001000010111011010101011011010110010000101101110; end
            14'd9735 : begin out <= 64'b0010101010010111101001101000110010011000011011101010101101010001; end
            14'd9736 : begin out <= 64'b0010011001111010001010011000001110101010101011101010001110011100; end
            14'd9737 : begin out <= 64'b1001110010100011000111101011011100101100000110010010010111001100; end
            14'd9738 : begin out <= 64'b0010100110010111100111110010111100101100001001100010000001101111; end
            14'd9739 : begin out <= 64'b0010010100100000001010100011011010100101111101010010100000011010; end
            14'd9740 : begin out <= 64'b0010101111000001001000100111000110001011101111100010001100100011; end
            14'd9741 : begin out <= 64'b1010100001001000001010100111010010101010101001001010110000000010; end
            14'd9742 : begin out <= 64'b0010011000000100001001011111000000101011010000001010011001010101; end
            14'd9743 : begin out <= 64'b1010101010000100100110001001001010101001101001111010101110010001; end
            14'd9744 : begin out <= 64'b0010000110000001101010110100001110100011110010011010000110000001; end
            14'd9745 : begin out <= 64'b0010010100000110101010110010000110101010111100111010100000000010; end
            14'd9746 : begin out <= 64'b0010010100101010001010010101001110100110001011110010011001110001; end
            14'd9747 : begin out <= 64'b1010011000001001100110000110100110100001101100011001000011100001; end
            14'd9748 : begin out <= 64'b0010100010001011001001000011101100100111100100011010000110001100; end
            14'd9749 : begin out <= 64'b1001110011101010000110101001011000101011000110010010100110110000; end
            14'd9750 : begin out <= 64'b1010101110111011101010110001000000100110000111001010101000010000; end
            14'd9751 : begin out <= 64'b0010001100010101101010100101100010100100100010001001100110101001; end
            14'd9752 : begin out <= 64'b1010100111000101101010001100111110101010110010101010010111101110; end
            14'd9753 : begin out <= 64'b0010101001001111001001001101000110100010001001000010101100010111; end
            14'd9754 : begin out <= 64'b0010010101010001101000001110100010101010101101011010100101100001; end
            14'd9755 : begin out <= 64'b0010011010100100101010000101100110101010001011001010011000101010; end
            14'd9756 : begin out <= 64'b0010101111111011001010000001111100100111001101110010010010001000; end
            14'd9757 : begin out <= 64'b1010011000011111001011000000110010100100101001000010100001110000; end
            14'd9758 : begin out <= 64'b0001110000111110001010100111000100101010111001111010011111010100; end
            14'd9759 : begin out <= 64'b0010001100000101001010010010111000100111101010100010001100000111; end
            14'd9760 : begin out <= 64'b0010011010100110101001000100011110101001000010010001110100100101; end
            14'd9761 : begin out <= 64'b0010100101000011100110110101000100100100110111010010000010011100; end
            14'd9762 : begin out <= 64'b1010100101110111001010011101011110101010000010110010011010000000; end
            14'd9763 : begin out <= 64'b0010110000010010001010111011011010101001101011111010010010001010; end
            14'd9764 : begin out <= 64'b0010010000010001101010000011011000100001011001110010010000110100; end
            14'd9765 : begin out <= 64'b0010011011001110001001101011001100101011101001101010100000110001; end
            14'd9766 : begin out <= 64'b1010011111000010001001111100000010100101111110101010010101101100; end
            14'd9767 : begin out <= 64'b1001110000110011101010011111001110101011010000101010100000011001; end
            14'd9768 : begin out <= 64'b1010100110011000001000100110001100101000101110111010101001111011; end
            14'd9769 : begin out <= 64'b0010010100101111000100011010001010101010001000011010101111010000; end
            14'd9770 : begin out <= 64'b1010100011000010001001111001000000101000101111010010011100110010; end
            14'd9771 : begin out <= 64'b1010011010011111001010101110011010101001111000001010101101100101; end
            14'd9772 : begin out <= 64'b0010001000001100101010111110001010100011100001101010101001110011; end
            14'd9773 : begin out <= 64'b1010101111001111101010011111100100100101000100000010010000111100; end
            14'd9774 : begin out <= 64'b1010100110100001101010111000010000100010011001100010010111000110; end
            14'd9775 : begin out <= 64'b0010100011010110101001111001111100011101111011101010011010111000; end
            14'd9776 : begin out <= 64'b1010010011100001001001110110000110101001101011110010010011100011; end
            14'd9777 : begin out <= 64'b0010010110010111101001001101101110101000011010000001000001000100; end
            14'd9778 : begin out <= 64'b0001111000000111001001011111101000011000110101011010010011001110; end
            14'd9779 : begin out <= 64'b0010100101011110101001000111101000101010001010111010101100111110; end
            14'd9780 : begin out <= 64'b1010101001011101101000111001101010101001101101010001110001110011; end
            14'd9781 : begin out <= 64'b0010100110111010001001001011001110010110110100011010100000101011; end
            14'd9782 : begin out <= 64'b0010011101101000001010011101001010100010010010011010011110001011; end
            14'd9783 : begin out <= 64'b0010010100001101101010000001011110101001000100100010100011110101; end
            14'd9784 : begin out <= 64'b1010010100100111001000110010001010101000100111001010100010101010; end
            14'd9785 : begin out <= 64'b0010101010011110101010111001001010101010011111010010101010000110; end
            14'd9786 : begin out <= 64'b0010101111010001001001000001011110011111010101110010011101011010; end
            14'd9787 : begin out <= 64'b1010010001000101101010011101100100101011011110100010100101101010; end
            14'd9788 : begin out <= 64'b0010011000001100101000111101001010100101001100010010010000111010; end
            14'd9789 : begin out <= 64'b1010101010110110101000100000100010101011010101011010100110100101; end
            14'd9790 : begin out <= 64'b0010100111000001001001001110000010101000000010110010101111111000; end
            14'd9791 : begin out <= 64'b0010011000011001001000000000110110100001011011000010100011010111; end
            14'd9792 : begin out <= 64'b0001111000000001101010111010101000101001000011101010101011111001; end
            14'd9793 : begin out <= 64'b0010101111100110001001111001010110101000011000110010011101100110; end
            14'd9794 : begin out <= 64'b0001010010110110001001111100000000100111001101110010100110010011; end
            14'd9795 : begin out <= 64'b0010011100001100000111001110000000101001110001111001111010101101; end
            14'd9796 : begin out <= 64'b0010101111110001000111000111011110100000001101110010000110111111; end
            14'd9797 : begin out <= 64'b1010101101110010101010111000010010100100001100001010010001001111; end
            14'd9798 : begin out <= 64'b1010001001011001100110101001111100001111010010001010010101101001; end
            14'd9799 : begin out <= 64'b1010100011000011101001101110110110101010111000110001110011011000; end
            14'd9800 : begin out <= 64'b1010100011111011001010110011001010010100111000000001101011111111; end
            14'd9801 : begin out <= 64'b0010101101100100101000110111101000101011010010001010000110100101; end
            14'd9802 : begin out <= 64'b0010001100001001101010110010110010101000101100000010011101110100; end
            14'd9803 : begin out <= 64'b1010101110110110101010011001101110101011111111110010101110011010; end
            14'd9804 : begin out <= 64'b1010101110111001101010100000100100011101011011011010100000001111; end
            14'd9805 : begin out <= 64'b1010101000110101001010100100010110100111011000101001001011110001; end
            14'd9806 : begin out <= 64'b0010100101100011100110000010100100100000111101100010100010100100; end
            14'd9807 : begin out <= 64'b0010100110000101001010100010011110101010111000000010100111110010; end
            14'd9808 : begin out <= 64'b0010100111000000101001111001100100100010011000011010101011001000; end
            14'd9809 : begin out <= 64'b0001011001001000101001000010011000100011001110110001111011000111; end
            14'd9810 : begin out <= 64'b1010011001010011101001100110101010100111110010000010011110110110; end
            14'd9811 : begin out <= 64'b1010100101100011001010110101110000100100101001010010100001100010; end
            14'd9812 : begin out <= 64'b1010100110010100101001011011010110101010111111001010000100001011; end
            14'd9813 : begin out <= 64'b1001101101010110101010101011011000011100100110000010001101100110; end
            14'd9814 : begin out <= 64'b0010100010101001000101011101000000100100011010100010011001101111; end
            14'd9815 : begin out <= 64'b0010101000111101001010101000110010101000001001100010101011111100; end
            14'd9816 : begin out <= 64'b1010100100001000001001111111001000100100010110000010101000111001; end
            14'd9817 : begin out <= 64'b1010100001100111001001011100010110101000011001010010010011100101; end
            14'd9818 : begin out <= 64'b1010101110110110000110011110000010101011011110000010101000101111; end
            14'd9819 : begin out <= 64'b0010100100001111101010100001000000100011110101001010001000111001; end
            14'd9820 : begin out <= 64'b0010101110111111101001000111110100101010101011000010100010110101; end
            14'd9821 : begin out <= 64'b1010011010001110001001101011011000100000010100011010100100111111; end
            14'd9822 : begin out <= 64'b1010100101111101101010000101011000101000110010010010011110111111; end
            14'd9823 : begin out <= 64'b1010011001111110001010110110001010000111001001001010100000101111; end
            14'd9824 : begin out <= 64'b1010011110101001101010000111010000011100100111000010100110110110; end
            14'd9825 : begin out <= 64'b0001110011000101101010111000110010101001100011101010000011111011; end
            14'd9826 : begin out <= 64'b1010101011111111101010011111000000101011011000001001101010010110; end
            14'd9827 : begin out <= 64'b0010011110000011101001011010001110100110011001100010100101000111; end
            14'd9828 : begin out <= 64'b1010101000111110101000101100101100100011011010100010011011011100; end
            14'd9829 : begin out <= 64'b1010010111001110101001011000111110100110000001011010100010010100; end
            14'd9830 : begin out <= 64'b1001110000101011001001101101100110100100000111110010010011011000; end
            14'd9831 : begin out <= 64'b1010001101001110101010010000000000100100001110010010101110100000; end
            14'd9832 : begin out <= 64'b0010011001111111100110001111101000101000101100000010010001101100; end
            14'd9833 : begin out <= 64'b1010101010000110100000000110011110101001001101000010100100010001; end
            14'd9834 : begin out <= 64'b0010011001001101000111010100100100100111010000111001110100100000; end
            14'd9835 : begin out <= 64'b1001011000110110000110011111010000011101100100001010101011100101; end
            14'd9836 : begin out <= 64'b0010101001010010100100110101010010100000000100001010010101110001; end
            14'd9837 : begin out <= 64'b1010101000100110001001001111001000100110101100000010010000010011; end
            14'd9838 : begin out <= 64'b0010011010111101101010101101001110100111001101111010001001000100; end
            14'd9839 : begin out <= 64'b1010100010000000001001100000101010101011101111001010001111001110; end
            14'd9840 : begin out <= 64'b0010110000010010001010100100010000101000100000100001110110111001; end
            14'd9841 : begin out <= 64'b1010011110100101101000110001100110100000001011011010101110101000; end
            14'd9842 : begin out <= 64'b0010010100000001101001011001011010011111000011110001110001111011; end
            14'd9843 : begin out <= 64'b1010100111001110101011000000100000101011011111111010011110011001; end
            14'd9844 : begin out <= 64'b1010010000111110101010101010111010011100010001000010010011011010; end
            14'd9845 : begin out <= 64'b0010100010100010101001011000001000100011101101101010011011010101; end
            14'd9846 : begin out <= 64'b0010010011011110001010001110110000101011110101001010101001011011; end
            14'd9847 : begin out <= 64'b0010011010111110101001100000110000101001100001100010010000110110; end
            14'd9848 : begin out <= 64'b0010101110011001101000000000100110101010100011100010100010011001; end
            14'd9849 : begin out <= 64'b0010101011101100001010010111001010101010011010110010010010000111; end
            14'd9850 : begin out <= 64'b1010110000001000001010111010100010100000100011101010101111110000; end
            14'd9851 : begin out <= 64'b0001110000110101101001110001011010101100001001000001111100011110; end
            14'd9852 : begin out <= 64'b0010010101101100001010001101001000101011011101100010101110110111; end
            14'd9853 : begin out <= 64'b1001100110011110101001100010011110100110100111000010101011100111; end
            14'd9854 : begin out <= 64'b0001010011110110001010000101011010101000000011001010010111001111; end
            14'd9855 : begin out <= 64'b0010000010011100101010001111111010010001100011101010100001000111; end
            14'd9856 : begin out <= 64'b0010100101000111001010100011000000101011001101001010010101111000; end
            14'd9857 : begin out <= 64'b0010110000111010101000010000110110100011001100011010011010011010; end
            14'd9858 : begin out <= 64'b0010100010011101001010100000000010101001011111010010000001001011; end
            14'd9859 : begin out <= 64'b0010000111000010101010010111001000101100010011101001001001101111; end
            14'd9860 : begin out <= 64'b1010101011001011100111111000001110101000101111101010100011111010; end
            14'd9861 : begin out <= 64'b0010000101000000101001010010110010101000110110111010010111101101; end
            14'd9862 : begin out <= 64'b0010100101001010001001111001101110101000111100001010101010000110; end
            14'd9863 : begin out <= 64'b0001100001110010000111100011110110101011000000010010010101101101; end
            14'd9864 : begin out <= 64'b1001111110000000101001111100101100101000010100101010010100100111; end
            14'd9865 : begin out <= 64'b0010101011010011101001000000111100101010001100000010000011100101; end
            14'd9866 : begin out <= 64'b1010100100110111101000001111010010101001010101110010101101111100; end
            14'd9867 : begin out <= 64'b0010011010000101101001000101101100101000001001000010101000011010; end
            14'd9868 : begin out <= 64'b1010101111010100001001011101000000100100000110100010100001110001; end
            14'd9869 : begin out <= 64'b1010011100111100001001001000111010100010001110101010011101011111; end
            14'd9870 : begin out <= 64'b0010010111110011001001011010010100100110001010010000000000101110; end
            14'd9871 : begin out <= 64'b1001110011101110101010111110000010100101000110000001100100010001; end
            14'd9872 : begin out <= 64'b1010010011001001001010000010110110101011010000110010101110001101; end
            14'd9873 : begin out <= 64'b0001111101110110001001011100001110101001100010101010101100000101; end
            14'd9874 : begin out <= 64'b1010101011001110101010111111110010100111010011000010011110110001; end
            14'd9875 : begin out <= 64'b1010101010101011100111101101010100100001100100101010100001010101; end
            14'd9876 : begin out <= 64'b1001111010001000100111111010001110101010001000011010100000110111; end
            14'd9877 : begin out <= 64'b1010000111110111101010110001101010100000000110011010011010110001; end
            14'd9878 : begin out <= 64'b0010100000001110101010001000111100101010000110001010101110011111; end
            14'd9879 : begin out <= 64'b0010011101110100101010000111110000100101111000101001111110101000; end
            14'd9880 : begin out <= 64'b1010101100010111001010100001001010101000000100100001111011101000; end
            14'd9881 : begin out <= 64'b0010001000110000101010001100110000011100010100100010000110110101; end
            14'd9882 : begin out <= 64'b0010100111110000101010101100101110100111111000011010100111001001; end
            14'd9883 : begin out <= 64'b1010100010011001001010111001000010011101001100100010101101000001; end
            14'd9884 : begin out <= 64'b1010101001100011001010110001011010100000010111001010011101101000; end
            14'd9885 : begin out <= 64'b1010010111111001000111010011100000011011010111000010100010010000; end
            14'd9886 : begin out <= 64'b1010101100001011001001011000001100101100010001010010001010011010; end
            14'd9887 : begin out <= 64'b0010100011100111101001011110111000011110111001011010000010100101; end
            14'd9888 : begin out <= 64'b1001101100011011100111000100111000100101111100110010010100001000; end
            14'd9889 : begin out <= 64'b1010011100100110101011000000001010100101000010010010101000000011; end
            14'd9890 : begin out <= 64'b0010010011011110001000010110110100101010100010011010100001110011; end
            14'd9891 : begin out <= 64'b0010101001001000001000111011010110101010110001001010001001010001; end
            14'd9892 : begin out <= 64'b0010100001011110101001101111011000101011010111000010101000110001; end
            14'd9893 : begin out <= 64'b1001100110101111000101110100001010011100010001100010000101110000; end
            14'd9894 : begin out <= 64'b0010100011100000100111001100000110101011101011011010011110111001; end
            14'd9895 : begin out <= 64'b1010011001000011001011000000001100011101100110010010101001101100; end
            14'd9896 : begin out <= 64'b1010000100111010101001000010000010100111111010100010100111001010; end
            14'd9897 : begin out <= 64'b0010100101100110001010011000101110101011100011100010101011100101; end
            14'd9898 : begin out <= 64'b1010100011100010001010101110101110011100110111111010000110000100; end
            14'd9899 : begin out <= 64'b0010101101000101101010110111001000011010100110110010101101000010; end
            14'd9900 : begin out <= 64'b0010101110101101001010100000011010011111110101101010100011010101; end
            14'd9901 : begin out <= 64'b1010000011001110001010000100101000101010100001111010101010011100; end
            14'd9902 : begin out <= 64'b0001101110100010101000010011011000101000010000000010010101001001; end
            14'd9903 : begin out <= 64'b0010101101101001001010011111000100101011000110000010100101000000; end
            14'd9904 : begin out <= 64'b1010000111010110001010010001101010100101000111101010011111111101; end
            14'd9905 : begin out <= 64'b1010101111110100001010101000000000101001000101110010100001010111; end
            14'd9906 : begin out <= 64'b0010101111011010001000001001101100101001011001001010011101111000; end
            14'd9907 : begin out <= 64'b0010100100011101101010110101111000101000110100010010100011100111; end
            14'd9908 : begin out <= 64'b1010011000010110100111011101000010100110000001100010101100100000; end
            14'd9909 : begin out <= 64'b0010100000111100001000011101000100101001000101011010101100111011; end
            14'd9910 : begin out <= 64'b0010010110110101001010110101011110101000000011011010100011100101; end
            14'd9911 : begin out <= 64'b1010100111010011000111110100110010100100110111101010011100001000; end
            14'd9912 : begin out <= 64'b1010101000010100001010010100111010011011001111001010011001001010; end
            14'd9913 : begin out <= 64'b1010010011110010101010110001001000101000101000011010110000011110; end
            14'd9914 : begin out <= 64'b1010010011110011101010011011010110100100000000011010010100000010; end
            14'd9915 : begin out <= 64'b0001111110001110101010001001001010101001100010111010101000000001; end
            14'd9916 : begin out <= 64'b1010100001111000001001010100101100101010011010101001001000010011; end
            14'd9917 : begin out <= 64'b0010100011001100001001110101010110101001001111101010100000101000; end
            14'd9918 : begin out <= 64'b1010101100111100101010010001010100000100010101111010100001101100; end
            14'd9919 : begin out <= 64'b0010100011011111101000101001101110100000011110000010000101001010; end
            14'd9920 : begin out <= 64'b0010001111101000001001011001011000101000101110100001111011000110; end
            14'd9921 : begin out <= 64'b0010010110011111100111010000111000101000011011111001101111001100; end
            14'd9922 : begin out <= 64'b0001000101001100001000001000110110101100000100100010100100001001; end
            14'd9923 : begin out <= 64'b0010000000100011101010000011000110100110100001011010011010010110; end
            14'd9924 : begin out <= 64'b1001111100111101000111001111100110010110111111011001110000011100; end
            14'd9925 : begin out <= 64'b1010100100101100001010111000110000100001000010111010011110000000; end
            14'd9926 : begin out <= 64'b1010101001010101101010000110111100101010101101011010100111011110; end
            14'd9927 : begin out <= 64'b0010101111010101101010011111001000100010011110000010101100111100; end
            14'd9928 : begin out <= 64'b1010101111011111101010010000111010101001101111001010100110110100; end
            14'd9929 : begin out <= 64'b0010101111000101001001011110010110101011011010100010101001101100; end
            14'd9930 : begin out <= 64'b0010100110110010101010101001011110101011100001011010101110011111; end
            14'd9931 : begin out <= 64'b0010101010011011001010111010111110101001101111101010001001111110; end
            14'd9932 : begin out <= 64'b0010100100100110001010011100000010100110000000011010100110101100; end
            14'd9933 : begin out <= 64'b1010100111011010001010101101010110100011100110111010101110111101; end
            14'd9934 : begin out <= 64'b0010101110010101101001001001101010101000001111001010010101000010; end
            14'd9935 : begin out <= 64'b0010101010001111001001100111010100101000000011110010101000111100; end
            14'd9936 : begin out <= 64'b1010100000001000001001101011000010100000101000011010100101111001; end
            14'd9937 : begin out <= 64'b0010101011110110001010001111100100101000010100001010010000010000; end
            14'd9938 : begin out <= 64'b1010010001001010001001010111111100101011010110100010100011001000; end
            14'd9939 : begin out <= 64'b0010101001000010000110110000111000101011011011010010011011011101; end
            14'd9940 : begin out <= 64'b1001101000100010101001101100011110100001011010000010010001100001; end
            14'd9941 : begin out <= 64'b1010001000000111001000000010101000011111100111110010101100001100; end
            14'd9942 : begin out <= 64'b0001010101000111101010111101111010011111011111110010101111001001; end
            14'd9943 : begin out <= 64'b1010000100100101001010111000000100101011000110000001110101101110; end
            14'd9944 : begin out <= 64'b1010101110001101001001011110001010101001100111111010001101001010; end
            14'd9945 : begin out <= 64'b1010100110111011100110110001000100101000111111011010011011011111; end
            14'd9946 : begin out <= 64'b0010011011111001101010101011111000101010011101110010010000010001; end
            14'd9947 : begin out <= 64'b1001101110001010101010101110110010100100111101010010100111101001; end
            14'd9948 : begin out <= 64'b0001101100010011101000101111000110101000001110101010100011100001; end
            14'd9949 : begin out <= 64'b1001111111011101001010111010111010100111111111110010100110000110; end
            14'd9950 : begin out <= 64'b0010101111000101001010001101010000101011101000111010100000010101; end
            14'd9951 : begin out <= 64'b1010010001111111101010010111101010100110111111010010000110110111; end
            14'd9952 : begin out <= 64'b1010001100011101001010001010101110100101001100011010100000101100; end
            14'd9953 : begin out <= 64'b1010100111010111101001111110001100100111011111011010101001010001; end
            14'd9954 : begin out <= 64'b0010101110010110101000001000011010010110001000101010100100001110; end
            14'd9955 : begin out <= 64'b0010100000011110101010111101101010100001100101101010100001011110; end
            14'd9956 : begin out <= 64'b0010011011000101101000111100101110100110001011101010101101011100; end
            14'd9957 : begin out <= 64'b1010101101100010000111010111011100100010010111110010010110011110; end
            14'd9958 : begin out <= 64'b1010010001110010101000101000010010101011010000110010000000110000; end
            14'd9959 : begin out <= 64'b1010000001010110001010011111011110100000011000011001110001001010; end
            14'd9960 : begin out <= 64'b1010000111010100001010011001001110011011100101010010010111111001; end
            14'd9961 : begin out <= 64'b1010001111010101100011011100111010100000010011111010101001110101; end
            14'd9962 : begin out <= 64'b1010001111011101001010100100101100101010111001111010100010000011; end
            14'd9963 : begin out <= 64'b0010100111101101100110111111110100100011110111101001110100001011; end
            14'd9964 : begin out <= 64'b0010100101100101101000100111011100100101100110110010101001111110; end
            14'd9965 : begin out <= 64'b0010001110010111101010001000010000011111111101111010101000111010; end
            14'd9966 : begin out <= 64'b1010100111110001101010001000000110101011110111001010100110000000; end
            14'd9967 : begin out <= 64'b1010000000001101101000000101111000101011110100001001110110100000; end
            14'd9968 : begin out <= 64'b0010100010010010101001000001010100100101011000000001101110000010; end
            14'd9969 : begin out <= 64'b0010010001111110101010010000101000101001001010110010100100100100; end
            14'd9970 : begin out <= 64'b0010100001010111001010111011010110101000000100110010011100011101; end
            14'd9971 : begin out <= 64'b1010001000011000101010110110110100100001010001111010100101111000; end
            14'd9972 : begin out <= 64'b1010010011001011101001011010010010101000010001100010000100010001; end
            14'd9973 : begin out <= 64'b1010101001001000100111111001010100101000100001110010000100100110; end
            14'd9974 : begin out <= 64'b1010110000010110001010011000100110101010001101111001101000101010; end
            14'd9975 : begin out <= 64'b0010000100110100101010100010100100101011111000000010011101111011; end
            14'd9976 : begin out <= 64'b0010101100001001000111001011101010101011110111111010100110101111; end
            14'd9977 : begin out <= 64'b1010010111110101101000110000110110100100001011111010100000010010; end
            14'd9978 : begin out <= 64'b1010101100111001101001011100111000101010101100011001011111011010; end
            14'd9979 : begin out <= 64'b0010010001100011001001000111001110101001100001010001000011100110; end
            14'd9980 : begin out <= 64'b1010101101101000001010001010110000001010110010010010011010110111; end
            14'd9981 : begin out <= 64'b1010101010010010101010010111000110100110110111111010010011001101; end
            14'd9982 : begin out <= 64'b0001011000100001001000110001110010010011110010111010010011001001; end
            14'd9983 : begin out <= 64'b1001110000100010101001000110110100101100000010000010100000001010; end
            14'd9984 : begin out <= 64'b0010100011111110001010010011010000100110100001011010101111111000; end
            14'd9985 : begin out <= 64'b0010101101001111001001011000110100101011101000111010100010001000; end
            14'd9986 : begin out <= 64'b0010101111011100101010011000110100101010001100010010101001011011; end
            14'd9987 : begin out <= 64'b1010001001001100101010000100101100101100011000101001110001011111; end
            14'd9988 : begin out <= 64'b0010100111000000001010100010000100101000111110001010100101001100; end
            14'd9989 : begin out <= 64'b0010100010010101001001011011001000100100010001011010011011100100; end
            14'd9990 : begin out <= 64'b0001110100101101100111000100111100101000101011000010100011000010; end
            14'd9991 : begin out <= 64'b1010100110101101101010110010100100100111101000001010011010111010; end
            14'd9992 : begin out <= 64'b0010001011111011101010010001101100100101100010010010100011000111; end
            14'd9993 : begin out <= 64'b0010101111010011001010100110011110101010011101101010100111110000; end
            14'd9994 : begin out <= 64'b1001111001101001001011000101010100101010001000000010101110010001; end
            14'd9995 : begin out <= 64'b1010100110100110101001100101110110101001000000010010100101101101; end
            14'd9996 : begin out <= 64'b0010101101000111101001010010110110101010111110001010101111011010; end
            14'd9997 : begin out <= 64'b1010101101000110001010100001010010101000010100010010101100000110; end
            14'd9998 : begin out <= 64'b1001101100110100001010111011110010100110001000100010011010101101; end
            14'd9999 : begin out <= 64'b0010011101111000001001110001001100101011001010111010011011010100; end
            14'd10000 : begin out <= 64'b1001100110000100001001010111000110100010100011101010001010101000; end
            14'd10001 : begin out <= 64'b1010010001000001001010000110010000100100011101010010100001110111; end
            14'd10002 : begin out <= 64'b0010101011101001001010100010001010101010001111010010100101001010; end
            14'd10003 : begin out <= 64'b0010100100010001000100111001000110101000001101100010011100010100; end
            14'd10004 : begin out <= 64'b1010001001100111001001100001101110101011100101101001110100111010; end
            14'd10005 : begin out <= 64'b1010100110001100001010100110100100100010001111001010011110011000; end
            14'd10006 : begin out <= 64'b1010100110111011101001000110111010100101110010001010100010101110; end
            14'd10007 : begin out <= 64'b1010101111111000001010101100011010101011011100111010001011101110; end
            14'd10008 : begin out <= 64'b0010001000100100001010101011000110100111001000000010010111111111; end
            14'd10009 : begin out <= 64'b0010010101100111101010010011010010101011010000111001100100100001; end
            14'd10010 : begin out <= 64'b0010100101000001101010110110111010101000100010000010000110100000; end
            14'd10011 : begin out <= 64'b0001111001001111001010011111100000101011000001001010011110001100; end
            14'd10012 : begin out <= 64'b1010010100101010001001110011110010101011001000111010101000011000; end
            14'd10013 : begin out <= 64'b1010100110010110101010000000100010100000001100100010101000010110; end
            14'd10014 : begin out <= 64'b1010011010010010000111010000011010011011100111110010101010101111; end
            14'd10015 : begin out <= 64'b0010100100011101101010101000111010100110101111000010100100101111; end
            14'd10016 : begin out <= 64'b1010000101101010101010100111010000101011111001110010100110110110; end
            14'd10017 : begin out <= 64'b1010101010000110001010010100110110011110010110101010101100001010; end
            14'd10018 : begin out <= 64'b0010101000010110001010010001110100101001100111111010010100000100; end
            14'd10019 : begin out <= 64'b1010101100110000100110111000010000101100010010000010011101100000; end
            14'd10020 : begin out <= 64'b1010010100100010001010000111011000101000001110110010011111011001; end
            14'd10021 : begin out <= 64'b0010010110110010101010001010010110100110100100000010101110010100; end
            14'd10022 : begin out <= 64'b1001100011101001101010010000101110011011011010100010101001110001; end
            14'd10023 : begin out <= 64'b0010000000000011101001001000001110101011011111010010100011011111; end
            14'd10024 : begin out <= 64'b1010100111100010001010101110101100101000011110101010100001001101; end
            14'd10025 : begin out <= 64'b0010101101100010001001001100000100101000100011101001110111011011; end
            14'd10026 : begin out <= 64'b0010011011110001001001010011010100101001100010001010001011100000; end
            14'd10027 : begin out <= 64'b1010100110010101001010010000010100101010000011111010000111110111; end
            14'd10028 : begin out <= 64'b0010100110000100001011000010101100100110001011110010010110010010; end
            14'd10029 : begin out <= 64'b0010101001101000001010100111001000010101010000001010100011001100; end
            14'd10030 : begin out <= 64'b0010100001001100101010011110001110101000111010001010001111001101; end
            14'd10031 : begin out <= 64'b1000111110001000101001010010111110100100111100110010011101110011; end
            14'd10032 : begin out <= 64'b1010010000111110001010010010000000100110001000111010000101100010; end
            14'd10033 : begin out <= 64'b0001100000000110001001011101101000101010100000110001111001000100; end
            14'd10034 : begin out <= 64'b1010101000011100101001111110011110101000010110000001101011000111; end
            14'd10035 : begin out <= 64'b1010011100000101101001010000001110011101000110011010100010010010; end
            14'd10036 : begin out <= 64'b1010101010010000001000001000111000101010011010111010101000011111; end
            14'd10037 : begin out <= 64'b1010101110111001101010100001100010101001110010011010101101100101; end
            14'd10038 : begin out <= 64'b0001100011110010100110100101101010101011000111000010010110110010; end
            14'd10039 : begin out <= 64'b1010010111100010001010001110000100011100011001001010101010001010; end
            14'd10040 : begin out <= 64'b0010010011100011100100110011001100100001111110101001111100000000; end
            14'd10041 : begin out <= 64'b1010011010101101000111001101101010100100100110010010001101000101; end
            14'd10042 : begin out <= 64'b1010010111110000000100100011111000100100100111101001110101001010; end
            14'd10043 : begin out <= 64'b1010001010110110001000011000111010101000111011011010000110000000; end
            14'd10044 : begin out <= 64'b0010000011111110001000011111010110101010011110000010100010110001; end
            14'd10045 : begin out <= 64'b0001111000101110101010111011001110101011000010010010101111101110; end
            14'd10046 : begin out <= 64'b0010011010011000101010000100100000101010011001001010101101111111; end
            14'd10047 : begin out <= 64'b0010100110000110101010001100111110101000101100101010000110100100; end
            14'd10048 : begin out <= 64'b1001100110101000101010011100111110100101101111111010101101101110; end
            14'd10049 : begin out <= 64'b0010100000110111001010100001001000101001011101000010001011111110; end
            14'd10050 : begin out <= 64'b0010100101101001001001111001101010100110100111010010010010111111; end
            14'd10051 : begin out <= 64'b0010011100111111101010101011111110101001111011101010100110100100; end
            14'd10052 : begin out <= 64'b0010101010111111101010011100010100101000011111101001110100100100; end
            14'd10053 : begin out <= 64'b0010100101101010001010110111101010101011100000000010101000000101; end
            14'd10054 : begin out <= 64'b1010101000010001101011000001001100101001111010101001110000011001; end
            14'd10055 : begin out <= 64'b0001100101111011001010110101000000101000111100000010101101111100; end
            14'd10056 : begin out <= 64'b1010100011100110101010000101111000011010110011101010000010110001; end
            14'd10057 : begin out <= 64'b0001101101000110001010000001001100101000001111110010010010011010; end
            14'd10058 : begin out <= 64'b1010001011001110001010001100101000100101010001011010100100011111; end
            14'd10059 : begin out <= 64'b1010010011000111101010100101010110101010110101111010001000000001; end
            14'd10060 : begin out <= 64'b0010100000100010101001010001110110010100111000010010000010001100; end
            14'd10061 : begin out <= 64'b0010011010001000101010110110001010101001001010011010101111001111; end
            14'd10062 : begin out <= 64'b1010011101011101101010111000001110100110011011000010011000110010; end
            14'd10063 : begin out <= 64'b0010100101011000000111110001011100101010000010111001110000000111; end
            14'd10064 : begin out <= 64'b0010101010111010001010001111000110100000100101110001110111011110; end
            14'd10065 : begin out <= 64'b0010101001011000101010100111011100100000010000001010101100000100; end
            14'd10066 : begin out <= 64'b1001111011000001101010110110000100101001101010010010001110010101; end
            14'd10067 : begin out <= 64'b0010011110000101100011101000011100100111100101001001011110100001; end
            14'd10068 : begin out <= 64'b1010101100101000100110100110000000100100101110101010011011010101; end
            14'd10069 : begin out <= 64'b0010100001110001101010101001011000100100101100101010011010010100; end
            14'd10070 : begin out <= 64'b1010101110110011001011000110001010100000100110001010101101010101; end
            14'd10071 : begin out <= 64'b1010010011000110001010000011111110101011000000111010000000100000; end
            14'd10072 : begin out <= 64'b0010101110111001001010110101111100011001111101111010001001110010; end
            14'd10073 : begin out <= 64'b0001100100011010001001110111101100101000110000001010100011100100; end
            14'd10074 : begin out <= 64'b0010101101101101101010110000000100101010101000110001111111100001; end
            14'd10075 : begin out <= 64'b0010101010011111101010101110111000101010010011100010011101100001; end
            14'd10076 : begin out <= 64'b1010101111100000001011000101100000101001111010000010100111001010; end
            14'd10077 : begin out <= 64'b0001010111001100000111100100100110100100100111100010100101001111; end
            14'd10078 : begin out <= 64'b1010101101110010101001111010011110101011011000010010101010101011; end
            14'd10079 : begin out <= 64'b1010010110001101101010000011110110101001001001001010011101100101; end
            14'd10080 : begin out <= 64'b0010010110110000001010101010011000101000100111000010101011111011; end
            14'd10081 : begin out <= 64'b1010101010010010101000001100110000100111000111010010101001101000; end
            14'd10082 : begin out <= 64'b1001101011000110101001101001100100101011100110101010011001011011; end
            14'd10083 : begin out <= 64'b1010101000001101001010100110011000100100001011011001000010011111; end
            14'd10084 : begin out <= 64'b0010101011011110001010100000101100100111010001111010101011101100; end
            14'd10085 : begin out <= 64'b0010100111110000101001111100000110011110000011100010010011010101; end
            14'd10086 : begin out <= 64'b0001110101111011101001001101011010100110011010001010001100001010; end
            14'd10087 : begin out <= 64'b1001110111101110101000011111110000101010100001101001101000100010; end
            14'd10088 : begin out <= 64'b0010100000000110001010011010101100101011000001101010100010101000; end
            14'd10089 : begin out <= 64'b1010100100101100101001111001111110100111011000001010011011110101; end
            14'd10090 : begin out <= 64'b0010101011000000000111100011010100101001100000011010010011101100; end
            14'd10091 : begin out <= 64'b1010100010001100101001111010111110101011000101101001100011100011; end
            14'd10092 : begin out <= 64'b1001111101101100100110110110000110101011101111111010010001000010; end
            14'd10093 : begin out <= 64'b0010101000100110101010000010100000101001110101011010100100000010; end
            14'd10094 : begin out <= 64'b1010100110010001001010111110111100011001111001001010101101100011; end
            14'd10095 : begin out <= 64'b0010011101001100100111011000101010101011001100110010011111100101; end
            14'd10096 : begin out <= 64'b1010100001000111001001011010111000011010000111110001001101110000; end
            14'd10097 : begin out <= 64'b0010101000000111001000110010011010101011100001111010001100100101; end
            14'd10098 : begin out <= 64'b1010010110001010001001100100000010100100000010011010100010100011; end
            14'd10099 : begin out <= 64'b1010100000011110101010000000001100101011101010110010001110000110; end
            14'd10100 : begin out <= 64'b0001111100111101101010011111000110100111011010110010011010000111; end
            14'd10101 : begin out <= 64'b1010010100000101001010001101000100101001011010101010011100100100; end
            14'd10102 : begin out <= 64'b0010101111101001001000100111110010101011111010011010100001010000; end
            14'd10103 : begin out <= 64'b1010010110101111001010111011110010100001101101101010100110000111; end
            14'd10104 : begin out <= 64'b0010101011100110001010100000100110011110011101001010001000110010; end
            14'd10105 : begin out <= 64'b0010101001100000001010000010001010100110000111010010010010010110; end
            14'd10106 : begin out <= 64'b1010000111111100101010000100110010010100010101011010001010010111; end
            14'd10107 : begin out <= 64'b0010100010111011001010000000000000010101111101000010101111111110; end
            14'd10108 : begin out <= 64'b1010100110010000101001111111010010101010101001101010101000111111; end
            14'd10109 : begin out <= 64'b0010100001001010101010101110011000100111100110110010001011111010; end
            14'd10110 : begin out <= 64'b0010001101111110101010100110010110101001010010001010101110100010; end
            14'd10111 : begin out <= 64'b0010101101111001001001010001011100101001100011011010100100011000; end
            14'd10112 : begin out <= 64'b1010000111101010001011000001111110101010011110001001111111111111; end
            14'd10113 : begin out <= 64'b0010010100000100001000101010100100100110011011010010010011111011; end
            14'd10114 : begin out <= 64'b0010100000000000001000100011001000101010000011110010000001111110; end
            14'd10115 : begin out <= 64'b1010100111111001100111000010111110100100111001101001110010011110; end
            14'd10116 : begin out <= 64'b0010010011010010001001000011110000100111011010111010101010011000; end
            14'd10117 : begin out <= 64'b0010011010111101100110001011001010100011010110010010100000111110; end
            14'd10118 : begin out <= 64'b1010000001001100100111011110100110010000001011001010001001001001; end
            14'd10119 : begin out <= 64'b1010001000010000001000100111001000100111001100011010101001000000; end
            14'd10120 : begin out <= 64'b0001100011111100101000111001010000100001001001110010100110110101; end
            14'd10121 : begin out <= 64'b1001110111110100001001111001100110101010101011011010000001001001; end
            14'd10122 : begin out <= 64'b0010001000111100101010101110100000101010101111100010100010110100; end
            14'd10123 : begin out <= 64'b0010010100101000100111101011111100101001001000110010101100100011; end
            14'd10124 : begin out <= 64'b1001111110100001101010110001111010101010111011001010011100101100; end
            14'd10125 : begin out <= 64'b1001011100001010001010101000000000101011011000101010101111101111; end
            14'd10126 : begin out <= 64'b1010011011001011101011000100101100100101100110011001111110001000; end
            14'd10127 : begin out <= 64'b0001011100011001101010101010100010101001001111101001110101010010; end
            14'd10128 : begin out <= 64'b1010010100110001101010010110100000100011101100101010001110011100; end
            14'd10129 : begin out <= 64'b1010011111000011000111001100001010100101000010010010100111110010; end
            14'd10130 : begin out <= 64'b0001111101100111100010110011010010100100011001011010010001111001; end
            14'd10131 : begin out <= 64'b0001111100111011101010110110101110100111100111110010010011000011; end
            14'd10132 : begin out <= 64'b0010100011100101100111101101010010101001100001110010100000110000; end
            14'd10133 : begin out <= 64'b0010011110011111001000110111110110101000000000100010011111111111; end
            14'd10134 : begin out <= 64'b1010100010110010101001010000010000100111111011011010101011101010; end
            14'd10135 : begin out <= 64'b1001111000110010001000110111010000101000011001100010101111000100; end
            14'd10136 : begin out <= 64'b0010010110000011001001111000010000100110000101001010101011011011; end
            14'd10137 : begin out <= 64'b1010100000100110101010000000100100101011010101110010100111010100; end
            14'd10138 : begin out <= 64'b1010100011000111001001100111110100101001110001111010100010100001; end
            14'd10139 : begin out <= 64'b0001111100100101001000010000001010101001010001001010101110100100; end
            14'd10140 : begin out <= 64'b0010100100111001001000011011001110100110110010111010100000000110; end
            14'd10141 : begin out <= 64'b0010101011101001001010001101101110101000010011010010101101001001; end
            14'd10142 : begin out <= 64'b1010101001011001100111010101100100101000001011010010010010000100; end
            14'd10143 : begin out <= 64'b0001111001110000101010000011110000100100110111000010101100011010; end
            14'd10144 : begin out <= 64'b1010100001001110101001011000001010101010100010011010010100001011; end
            14'd10145 : begin out <= 64'b1010101011111100001010010011000010100011110010100001110101010111; end
            14'd10146 : begin out <= 64'b1010001001110110000100101001101110010101011000001010101000010000; end
            14'd10147 : begin out <= 64'b1010001110110111101001111101011100101001010101010010101010011100; end
            14'd10148 : begin out <= 64'b1010100101011000001010001100101000010011010111011010101100110010; end
            14'd10149 : begin out <= 64'b1010100101000010001010011001010110100101000000000010011010100111; end
            14'd10150 : begin out <= 64'b0010100001000111001010110001110110011101000111010010100011111111; end
            14'd10151 : begin out <= 64'b0010100100110001100111011000000010101010111011101010101111011110; end
            14'd10152 : begin out <= 64'b0010010101001110101010010100010000100101101010111001111100111011; end
            14'd10153 : begin out <= 64'b1010100011000111101010010100101100100110000110000010011100010011; end
            14'd10154 : begin out <= 64'b0010010001111000100111100001110000100100000101001010000001100110; end
            14'd10155 : begin out <= 64'b0010100001110010001010100100011110100101000101011010101100101001; end
            14'd10156 : begin out <= 64'b1010100110110101101001010011100100100100010110011010100011100111; end
            14'd10157 : begin out <= 64'b0010101111110000101001101100100000100100100000000010100011100011; end
            14'd10158 : begin out <= 64'b0010100000110001101001001100000010101010000011001010100011110000; end
            14'd10159 : begin out <= 64'b0010100101110011000101111001111100100010100101110010101111001001; end
            14'd10160 : begin out <= 64'b0010101100100010001001011001001110101011010010001010010111100011; end
            14'd10161 : begin out <= 64'b1010101110110101101010010110011110101000111011001010010101101110; end
            14'd10162 : begin out <= 64'b1010101010110101101000010010101100101010111001111010011110011100; end
            14'd10163 : begin out <= 64'b0010101111110010101011000001101100100000011011100010011110011100; end
            14'd10164 : begin out <= 64'b0010011000011101101010000110001110101001111111100010000100111111; end
            14'd10165 : begin out <= 64'b1010011000011101101000010000000000100010110111101010001001011000; end
            14'd10166 : begin out <= 64'b1010011101001100101000110001100110100110000001100010101001010011; end
            14'd10167 : begin out <= 64'b0010011100111001101010001100001010101011011001000010011111100110; end
            14'd10168 : begin out <= 64'b0010010111001111001001110101110100101000100000100001111100000010; end
            14'd10169 : begin out <= 64'b1010010111001000101001100011010000101011000110111010000101001110; end
            14'd10170 : begin out <= 64'b1010011111101100100100010000011000101001001110110010100011010101; end
            14'd10171 : begin out <= 64'b1010100111101010101010100101101100101011111000000010100111010011; end
            14'd10172 : begin out <= 64'b0001010100011010001010000010001010101001011000000010000010110000; end
            14'd10173 : begin out <= 64'b1010101000010010101001010000010100100101010011000010100000100001; end
            14'd10174 : begin out <= 64'b1010101000001011001010001111101000101001011110000001111111111011; end
            14'd10175 : begin out <= 64'b0001110101101111101010011011011000100111001101110001111101111001; end
            14'd10176 : begin out <= 64'b0010101100100101101010101110000110101010010010000010101110011100; end
            14'd10177 : begin out <= 64'b1010011111111101001001011111110000101011000111100010101100101010; end
            14'd10178 : begin out <= 64'b0001010011101000000111100100111110100101011101110010100011010110; end
            14'd10179 : begin out <= 64'b0010001100100001101001000110110010100111000011111010001101110111; end
            14'd10180 : begin out <= 64'b0001110010000010001010111011010100100100101111011010100011001100; end
            14'd10181 : begin out <= 64'b1010100111101101001010100111100110101001101111110001110010101001; end
            14'd10182 : begin out <= 64'b1010101110010011101001110110010110101011100000010010101000001011; end
            14'd10183 : begin out <= 64'b1010010100110011101010001111100010101011001110010010011111100111; end
            14'd10184 : begin out <= 64'b1010011001011100001001010110111010011111110111011001101100010100; end
            14'd10185 : begin out <= 64'b1010000000010010101001011100100110101000100100010001100100101100; end
            14'd10186 : begin out <= 64'b0010101010110101101010110110111010011110101101100001000000000100; end
            14'd10187 : begin out <= 64'b1010001000110000001000111100100000100010001111011001010011010110; end
            14'd10188 : begin out <= 64'b1010011110010011101001000100011110011110111011100010100110011101; end
            14'd10189 : begin out <= 64'b1001001101010110001010111110110110101011001100111010001111110101; end
            14'd10190 : begin out <= 64'b1010101011000110100101010110001000101010000100111010011101010111; end
            14'd10191 : begin out <= 64'b0010100110010000001010010111110010101011010000001010101011110000; end
            14'd10192 : begin out <= 64'b1001001110011000001010010000011000101001110011111010000011000110; end
            14'd10193 : begin out <= 64'b0010100011100101101001100110110010101010100011001010011101010010; end
            14'd10194 : begin out <= 64'b1010101011001001001011000001110010100100100010000010010100000110; end
            14'd10195 : begin out <= 64'b1010100100111001001010000000100110101001100000111001111100100000; end
            14'd10196 : begin out <= 64'b1001100101010111001001110011010010101000000101001010100001101010; end
            14'd10197 : begin out <= 64'b0010000010100111001011000011100000101011001001011010011110011001; end
            14'd10198 : begin out <= 64'b1001111111001010001010100010101010100000011100110010001100011111; end
            14'd10199 : begin out <= 64'b1010011001011101001010000000101000100010000111000010101000000000; end
            14'd10200 : begin out <= 64'b0010101010110010001001000101010110101000110100110010010001110011; end
            14'd10201 : begin out <= 64'b0010101101000111001010101011111110101001011110101010100010110111; end
            14'd10202 : begin out <= 64'b0010101101111110101000101101010110101011000101100010101111010011; end
            14'd10203 : begin out <= 64'b1010101001010001101001000000010110101010001011100010100001010100; end
            14'd10204 : begin out <= 64'b0010100111011111101010000100100010100110110111000010001101110000; end
            14'd10205 : begin out <= 64'b0010101100100011101010101101010000101001010001011001011011000101; end
            14'd10206 : begin out <= 64'b1010100100011100101010011110000010100000101011110010000000010111; end
            14'd10207 : begin out <= 64'b0010000010101011101001111010111100101010100110000010011001001010; end
            14'd10208 : begin out <= 64'b1010101000101101001010101010011100101000100100100010101011010001; end
            14'd10209 : begin out <= 64'b0010011101011000001010101101111110100010010001011010101110010001; end
            14'd10210 : begin out <= 64'b1010011111011010001001100001000000100110110010001010001000110011; end
            14'd10211 : begin out <= 64'b1010100111000100101001111111110010101000001110110010011100011000; end
            14'd10212 : begin out <= 64'b0010010101111010101010010100110000101010001011100010101110010001; end
            14'd10213 : begin out <= 64'b1010000110110001001010011100011100101000010111011010011011011101; end
            14'd10214 : begin out <= 64'b1010010100000001001010111001100110100001110111100010010100110111; end
            14'd10215 : begin out <= 64'b0010100000111101101001001101011110100101000110100010101010011000; end
            14'd10216 : begin out <= 64'b1010100011001000101010000011100110011111010111111010010111111111; end
            14'd10217 : begin out <= 64'b0010011111101110001000000001000000101001000111010010001110000100; end
            14'd10218 : begin out <= 64'b0010100000000011100110111111010100100100010110011010010110101100; end
            14'd10219 : begin out <= 64'b0001101001001001100110000100011100101010011110000010100101000010; end
            14'd10220 : begin out <= 64'b1001011110110110001010010110110000100110110101111010011011101001; end
            14'd10221 : begin out <= 64'b0001111001010000101010011110010110101011110110010010101110000000; end
            14'd10222 : begin out <= 64'b0010100111001110101001010101101100100010100100101010101111110001; end
            14'd10223 : begin out <= 64'b0010000011010100101010101001001010101010011011001010011111011010; end
            14'd10224 : begin out <= 64'b1010001101110100001001000110011010100010101001001010010000001010; end
            14'd10225 : begin out <= 64'b1001110100011000101010001100000010100111011100011010100000101110; end
            14'd10226 : begin out <= 64'b0010000000110011101000010111001000100100000110111001100011000000; end
            14'd10227 : begin out <= 64'b0010100111000100101010011000110110101001110100000010001001111001; end
            14'd10228 : begin out <= 64'b0010001010101111101000101101100010100000001001110010101010001011; end
            14'd10229 : begin out <= 64'b1010100110110111101001000101001000101011110010011010011011000011; end
            14'd10230 : begin out <= 64'b1010010010011101101001001001101010101001001001111010010010011100; end
            14'd10231 : begin out <= 64'b1010100010100011001001000111111110100011110011001010100011011101; end
            14'd10232 : begin out <= 64'b1010101000010101101001111100011000010111110010001010101000110110; end
            14'd10233 : begin out <= 64'b0010100010000010101001001110001110101000101001011010001100100101; end
            14'd10234 : begin out <= 64'b0010101011100111101001100100001110100011100010001010100001001001; end
            14'd10235 : begin out <= 64'b0010100000101000000111110101010100101010001110011010011110010000; end
            14'd10236 : begin out <= 64'b0010100101100011101010101100001010100111101111100010100100001100; end
            14'd10237 : begin out <= 64'b0010100011011001101010111010010010100100111000011010101011111101; end
            14'd10238 : begin out <= 64'b1010101011100011101001010101001000101000001111011010010110011111; end
            14'd10239 : begin out <= 64'b0010100001111110001010001001101010100101000111011010011011000111; end
            14'd10240 : begin out <= 64'b0010101011110001001000110101100000100100001111111010000111110011; end
            14'd10241 : begin out <= 64'b0010001110110010001001101100010000101000100010100010100001011101; end
            14'd10242 : begin out <= 64'b0001101100110101101010100001101110101001111100000010010110000110; end
            14'd10243 : begin out <= 64'b0010101000110111001010101001011100001110011110010010100101001011; end
            14'd10244 : begin out <= 64'b0010001100111101101010011000111010101010111111100010100100000100; end
            14'd10245 : begin out <= 64'b1010000101011101100110001000010010011100001101101010010001110111; end
            14'd10246 : begin out <= 64'b1010101111110001101010000011110110101011110110010010011100001001; end
            14'd10247 : begin out <= 64'b1010101110110011001010110000011010101001000011101010001100110100; end
            14'd10248 : begin out <= 64'b0010000000011011101010000111000000101001001000000010100110101011; end
            14'd10249 : begin out <= 64'b0010100001100000101001100011010010101000000110011010010000101011; end
            14'd10250 : begin out <= 64'b0010010110011111001010110111110110100111001111100010010111110001; end
            14'd10251 : begin out <= 64'b1010100111101011001010101101010010100000010001000010101010110110; end
            14'd10252 : begin out <= 64'b0010011000101100001010010100011000101000001000010010101101101001; end
            14'd10253 : begin out <= 64'b0001111100010110001001011010111000100110000100111010101111101110; end
            14'd10254 : begin out <= 64'b1010100110100100001010111101000010101010001110100010100001110010; end
            14'd10255 : begin out <= 64'b1010011010110010101010101011110110101001001011101001110111110011; end
            14'd10256 : begin out <= 64'b0010010110010010100001010100000110101011101110110010100001010001; end
            14'd10257 : begin out <= 64'b0010100101101010101001000100000100101001110010110010101000001110; end
            14'd10258 : begin out <= 64'b1010101011000111101010111101001000100100101000111010000101000110; end
            14'd10259 : begin out <= 64'b0010011001011010101000010101011110101011110101111001011001001111; end
            14'd10260 : begin out <= 64'b0001110000111100001010100100100010101001000010111010011111010001; end
            14'd10261 : begin out <= 64'b0010010001100000001010000110111000011011011101110010101011110100; end
            14'd10262 : begin out <= 64'b1010100011110110001010110101110000101000001000011010100011100110; end
            14'd10263 : begin out <= 64'b0010101011011111101001001000011000100111001000111010100100100111; end
            14'd10264 : begin out <= 64'b1001110001101011001010110000110000100001111011010010100111100011; end
            14'd10265 : begin out <= 64'b1001011101010010001001011010011010101000011001111010100001100011; end
            14'd10266 : begin out <= 64'b1010010101110101101000000110101110100010110101011010100101110000; end
            14'd10267 : begin out <= 64'b1010100011000011001001100001010000101010001100000001110001000111; end
            14'd10268 : begin out <= 64'b1010000101010010001001010100101010011000110100101010100011010111; end
            14'd10269 : begin out <= 64'b1010011111000110001000011110011100100110111101101010101000000101; end
            14'd10270 : begin out <= 64'b1010100001000010001010010100010100101100011011000010101101001101; end
            14'd10271 : begin out <= 64'b0001110111000000001000100000011010101000101101111010100001100110; end
            14'd10272 : begin out <= 64'b1001100101111001101010010010111010100010100011010010001110001100; end
            14'd10273 : begin out <= 64'b1010101101100000101010000100001100101010010001110010101000101001; end
            14'd10274 : begin out <= 64'b1000101010000000001010000000100000101010111011010010100000111110; end
            14'd10275 : begin out <= 64'b0010000110010011101000011111111000101011001011011001111111101111; end
            14'd10276 : begin out <= 64'b0010011010100011001010100011011110101000011011000001111111111111; end
            14'd10277 : begin out <= 64'b1001110101001101001001010111000000100100101001010010101000111100; end
            14'd10278 : begin out <= 64'b0010100010001000001001111001100100100111101001101010100000000001; end
            14'd10279 : begin out <= 64'b1010100111101010001000100001111010101010011010111010100010110110; end
            14'd10280 : begin out <= 64'b1010100010111001101000110011010000101001010011101010100011010010; end
            14'd10281 : begin out <= 64'b1010100010000001101010101101101110100101100100100001110100001000; end
            14'd10282 : begin out <= 64'b0001101110111001101000111110000010101010011110001001111011100011; end
            14'd10283 : begin out <= 64'b1010101001110100001010101000011010100101111101111010011000111110; end
            14'd10284 : begin out <= 64'b1010010100001100001010000100100010011000111011111010011010111101; end
            14'd10285 : begin out <= 64'b1010000001110100001010101111100100100011000001101010100001111111; end
            14'd10286 : begin out <= 64'b1001111111110011001001100000010100100100001000010010100100011010; end
            14'd10287 : begin out <= 64'b0010101000001001001010001010001000101000000111000010011111101101; end
            14'd10288 : begin out <= 64'b0010101011001110001000011001100010101011000110010010010001100100; end
            14'd10289 : begin out <= 64'b0010101000111001101000100011001010101010111111001001111110111100; end
            14'd10290 : begin out <= 64'b0010001010011110001010110110011000100111100100110010101101011010; end
            14'd10291 : begin out <= 64'b1001101000111110101010101100011010101000000110001010010110011001; end
            14'd10292 : begin out <= 64'b0010001110010000101001000100111100011111110000000010101100100010; end
            14'd10293 : begin out <= 64'b1010011000111111001000100011001110101001001001110010010100011110; end
            14'd10294 : begin out <= 64'b1010101000111000101010111001110010101010100111100010100110100111; end
            14'd10295 : begin out <= 64'b1010010001010111001001100101110110100101100000000010011101101001; end
            14'd10296 : begin out <= 64'b0010101000101110101010110010101110101010111001100010101100011001; end
            14'd10297 : begin out <= 64'b1010011111010111101010001100010110101010010101011010100101101101; end
            14'd10298 : begin out <= 64'b1010011001010010001010000101101000100011011101011010000111010100; end
            14'd10299 : begin out <= 64'b0010100101100000101001001101000000101011000101001010100010000000; end
            14'd10300 : begin out <= 64'b0010010110101111101010001011000000100100110001001010101000110111; end
            14'd10301 : begin out <= 64'b1010010100010010000110101110111000101001010100011010011001000010; end
            14'd10302 : begin out <= 64'b0010010110110010101001011101100110011011011111000010011101001011; end
            14'd10303 : begin out <= 64'b0010000001110000101010001001001010101011010101100010011101001001; end
            14'd10304 : begin out <= 64'b1010010110001010100111101011110000101010000100110010101110110110; end
            14'd10305 : begin out <= 64'b1010001011000011101001000111010000100110100101111010100011111001; end
            14'd10306 : begin out <= 64'b1010100001111110101010011110100000101000011110010010100100000110; end
            14'd10307 : begin out <= 64'b1010101010010011101010001000011100101000011110101010010010110100; end
            14'd10308 : begin out <= 64'b1001111110001101101010110101111110100001101111111001001101010110; end
            14'd10309 : begin out <= 64'b1010100100100000101001010010011000100100000111010010101110001001; end
            14'd10310 : begin out <= 64'b0010011001101110101010011111000010101011011111000010100001100001; end
            14'd10311 : begin out <= 64'b0010101000001101001000000111001110100100111000010010100110010110; end
            14'd10312 : begin out <= 64'b1010100011101101001010111110001010100111110000110000001011000011; end
            14'd10313 : begin out <= 64'b0010110000001011101001001111100010100101010011000010011101110101; end
            14'd10314 : begin out <= 64'b1001110011000111001010010011000100011000010001100010101010001011; end
            14'd10315 : begin out <= 64'b0010010000101110001010010101110000101001110011101010101001110011; end
            14'd10316 : begin out <= 64'b0010100110100011001010111011001100100011000000001010100000110101; end
            14'd10317 : begin out <= 64'b1010100111001010101010100001001110101001001111000010100100100111; end
            14'd10318 : begin out <= 64'b1010101011010010001010001111011000011001100100000010011100001010; end
            14'd10319 : begin out <= 64'b1010100010101101001001000001101010100101111110111010100010000101; end
            14'd10320 : begin out <= 64'b1010101101100100001001111111011010101010000110111010101101000111; end
            14'd10321 : begin out <= 64'b0010100000000111001010010111010110100111000001100010101011010000; end
            14'd10322 : begin out <= 64'b0010100101010101001000111100000000101011001100101010000101110111; end
            14'd10323 : begin out <= 64'b1001101101011110101000000101100000100001110101101010101011000001; end
            14'd10324 : begin out <= 64'b1001110100100101001010111101011010101011100100111010101011010010; end
            14'd10325 : begin out <= 64'b0010001110110100101000001011101100100111100111111010100011000000; end
            14'd10326 : begin out <= 64'b0010011111101111100101111011010100101000100011100010011111000101; end
            14'd10327 : begin out <= 64'b0010100101010101001010101101001010101000100010111001111110010100; end
            14'd10328 : begin out <= 64'b0001110101110000101010111100110100101001100000100010011101100101; end
            14'd10329 : begin out <= 64'b0010000101010000001001001000000100101001010001010010100110111010; end
            14'd10330 : begin out <= 64'b1010101111100000101010100001000110101011001111110010010000010011; end
            14'd10331 : begin out <= 64'b1010100100110101000110111100110110011100111001101010101001011001; end
            14'd10332 : begin out <= 64'b0010101101100111001001100001101110101010000110100010101000101010; end
            14'd10333 : begin out <= 64'b0010100101000011001010011110111110101001110001101010101000111010; end
            14'd10334 : begin out <= 64'b0001111111111011001010011111110100101011100001001010101100100100; end
            14'd10335 : begin out <= 64'b1010100011000101001001001000111100101011111000101010010101101100; end
            14'd10336 : begin out <= 64'b0010010100101101100100010000111100101011110110110010101011011111; end
            14'd10337 : begin out <= 64'b1010100001100000001001011101011100100110101101110010100010110100; end
            14'd10338 : begin out <= 64'b0010100011011010001001011100111100011100010001010010101111100011; end
            14'd10339 : begin out <= 64'b0010000010001100101010111100111010101001110001110010101110011011; end
            14'd10340 : begin out <= 64'b1010011000011010001010001110011000011100111011100010011111111001; end
            14'd10341 : begin out <= 64'b1001101011001100101010100101010010101000100011001010010100101011; end
            14'd10342 : begin out <= 64'b0001110000001011101000101000010110010101111001001010100001001010; end
            14'd10343 : begin out <= 64'b1001100001110100001000010101011000101000001110001010001100001011; end
            14'd10344 : begin out <= 64'b1010101100110110101001000010111100101001100110000010000101011011; end
            14'd10345 : begin out <= 64'b1010100111100010101001100100101110101011000001101010100101010010; end
            14'd10346 : begin out <= 64'b0010010001100011001010001111110010101001000001000010011101110110; end
            14'd10347 : begin out <= 64'b0001101001010011101010001110101010100110000111101001111101011100; end
            14'd10348 : begin out <= 64'b1010101000100100000111111110011100100000111100111010101011001000; end
            14'd10349 : begin out <= 64'b0010011110000001101010010101110000101010110110001010100000100110; end
            14'd10350 : begin out <= 64'b0010011110101010001010100001101010100011001011111010100111011011; end
            14'd10351 : begin out <= 64'b0010011100011111100111011110001010100101011101110010000100101010; end
            14'd10352 : begin out <= 64'b0010011010111000101010000000011100100111000111000010100101010100; end
            14'd10353 : begin out <= 64'b1010010111011001100111000100001000100111101111001010010000101000; end
            14'd10354 : begin out <= 64'b0010100000110000101000010001101000010111001111000001111000110000; end
            14'd10355 : begin out <= 64'b0010100111001101101010111001010100100110010100100010100111000101; end
            14'd10356 : begin out <= 64'b1010001011100010001010011010001100100110011011100010010100110001; end
            14'd10357 : begin out <= 64'b0010000110110000001001011011100100100110100010110010100100100110; end
            14'd10358 : begin out <= 64'b1010101110110101100110011001010100100110100000010001111010101100; end
            14'd10359 : begin out <= 64'b1010101000011001001000111111000100101000100010100010110000111100; end
            14'd10360 : begin out <= 64'b0010011110011111001010010011101010101011011011000010101100001001; end
            14'd10361 : begin out <= 64'b0010000100111101101001101100100110101011001010101010011000010101; end
            14'd10362 : begin out <= 64'b1010100101001010001010011101000110100001001100101010011010110000; end
            14'd10363 : begin out <= 64'b0001010101010111101010100000101100100011111111100010100100111001; end
            14'd10364 : begin out <= 64'b1010011010111010001000000111101010101010010011000010101010111101; end
            14'd10365 : begin out <= 64'b1010100100011011001000000000110010100111101001101010100000101111; end
            14'd10366 : begin out <= 64'b1010101101000011101010010000001000100100011011001010010000101000; end
            14'd10367 : begin out <= 64'b1010100111000111101010111110001110100010001001111010100011101100; end
            14'd10368 : begin out <= 64'b0010001110110001101000010101101100101010110111100010100000111111; end
            14'd10369 : begin out <= 64'b0010010001010110001010011010010110100100111101010010100111100110; end
            14'd10370 : begin out <= 64'b1001100001010001100110111010000100100010010100110010101001101110; end
            14'd10371 : begin out <= 64'b0010101100111110101010111000100100100001000110011001110110001001; end
            14'd10372 : begin out <= 64'b0010101001011000001010110000110010011000101000000010011101010111; end
            14'd10373 : begin out <= 64'b1010010011001010100110111100010110101010011111000001010011111001; end
            14'd10374 : begin out <= 64'b1010010000100010000111100100001010100101001011010010100111101011; end
            14'd10375 : begin out <= 64'b0010100110100101101010001010011100101011100110010001111000100110; end
            14'd10376 : begin out <= 64'b1010101100111100001010110001100000101010111010110001010111100100; end
            14'd10377 : begin out <= 64'b0010010111001101100101010101111110101001111101010010010010000101; end
            14'd10378 : begin out <= 64'b0010010111110001001010010100000010010010101001010010101010101010; end
            14'd10379 : begin out <= 64'b0010011110010111101010011000000110101001101101010010100000000010; end
            14'd10380 : begin out <= 64'b0010100010111010101010010010100010101011010010110010001011111110; end
            14'd10381 : begin out <= 64'b0010100000111010001001110110110010101000110110010010100100111010; end
            14'd10382 : begin out <= 64'b0010010001100110100111000101000110101001100100110010010111001001; end
            14'd10383 : begin out <= 64'b1010100001101011101010110100001000101011000011100010010111101100; end
            14'd10384 : begin out <= 64'b1001111001110011101010011101111100101001110111111010101010110000; end
            14'd10385 : begin out <= 64'b1001100001101000001010100100111010101001110100011010101101011100; end
            14'd10386 : begin out <= 64'b1010100001100001101000100110001100100101110101011010101101001101; end
            14'd10387 : begin out <= 64'b0010101100100111101000010110110000101001011010011010101111100111; end
            14'd10388 : begin out <= 64'b1010100011010010001010011101101100101011100101111010101111010111; end
            14'd10389 : begin out <= 64'b0010011010011110101001101110000000101011001001101010000100101110; end
            14'd10390 : begin out <= 64'b0001101110100110101010100110010110011010110010000001111001110001; end
            14'd10391 : begin out <= 64'b1001101101010010101010110001010100101000110100110010101000110000; end
            14'd10392 : begin out <= 64'b0010011101101011100011010001001000101001100101000010000100101000; end
            14'd10393 : begin out <= 64'b0010100010011011001010011011101110101000111111011010001111001111; end
            14'd10394 : begin out <= 64'b1010011010101011101010101110110010011000100111000001111001101110; end
            14'd10395 : begin out <= 64'b1010001001100001101010010101110110101001100000011010010011110111; end
            14'd10396 : begin out <= 64'b1010010100001110101000110011011010101001111100001001101100100000; end
            14'd10397 : begin out <= 64'b1010100010000110001010010000000100011100001101010010100101000111; end
            14'd10398 : begin out <= 64'b1010001101011011101001110011110100100000100100011010001101111100; end
            14'd10399 : begin out <= 64'b1010101011110110101010000011101100100000110011100010100000000101; end
            14'd10400 : begin out <= 64'b0001101100110111101010110100101100100000101100110010010011100111; end
            14'd10401 : begin out <= 64'b0010001011000111001010011111100100100101111101000010010110111111; end
            14'd10402 : begin out <= 64'b1010001010101111001010100011000100101001010010001010101101010011; end
            14'd10403 : begin out <= 64'b0001111101111111001010011100011100100000001100001001011111110010; end
            14'd10404 : begin out <= 64'b1010100011111001101001111011111010101100000101011010010010000100; end
            14'd10405 : begin out <= 64'b0010001011010111101001011000010000101000011111000010010100000010; end
            14'd10406 : begin out <= 64'b0010010000111100001010010111000000101011001001000010010110110101; end
            14'd10407 : begin out <= 64'b0000110001001100101001101001111100100110010011111010101111011110; end
            14'd10408 : begin out <= 64'b1001010111011000001001010100000110101011001110100010011110010001; end
            14'd10409 : begin out <= 64'b1010100101001011101000101111001100100101110111010001111010101111; end
            14'd10410 : begin out <= 64'b1010100100101100101010010011110010101100000010100010101000111000; end
            14'd10411 : begin out <= 64'b0010010010000100101010111000101110101010111011110010000111010010; end
            14'd10412 : begin out <= 64'b0001100111100000101001110000010000100110001011000010010100001101; end
            14'd10413 : begin out <= 64'b0010100101000100100111111010011110100111100110001010011100000010; end
            14'd10414 : begin out <= 64'b0010011000110101001010101100101110100111010111100010100100011010; end
            14'd10415 : begin out <= 64'b1010100110110011101000111001111100101000001100101010100100111110; end
            14'd10416 : begin out <= 64'b1010011010000100001001110001011000100111110000100001011100001011; end
            14'd10417 : begin out <= 64'b1010000100111110101001100010011110101010011101001001110110011000; end
            14'd10418 : begin out <= 64'b0001010100110111000111100111011110101010001111000010000101011011; end
            14'd10419 : begin out <= 64'b0010101011101111001000100000011000101000000010001010101100011000; end
            14'd10420 : begin out <= 64'b1010101100110001101001101001001110100100110110111010011001110011; end
            14'd10421 : begin out <= 64'b1001101100000111101010110000110010101011110110101010101110011101; end
            14'd10422 : begin out <= 64'b0010101000001010101010010011111100101011000101011010000111110101; end
            14'd10423 : begin out <= 64'b0010101000111110001001011000011000101010110111100010011100011010; end
            14'd10424 : begin out <= 64'b1001010001100011101010011010101010101011110000001010100010011101; end
            14'd10425 : begin out <= 64'b0010101101110111101010000100101010100101001101011010000111011110; end
            14'd10426 : begin out <= 64'b1010101001110110101010101110001010100011010100100010100010101101; end
            14'd10427 : begin out <= 64'b1010100011010111001010001110100100101001011100101001010001101000; end
            14'd10428 : begin out <= 64'b1010100111101001001010101001011000101010101111001010100010010010; end
            14'd10429 : begin out <= 64'b1010100001111010001010111110000000101011001101000010101001110101; end
            14'd10430 : begin out <= 64'b1001111101001101101010000011100110101100000000010010010001011011; end
            14'd10431 : begin out <= 64'b0010010100100010000110100001110110101000010110011010000011111001; end
            14'd10432 : begin out <= 64'b0010110000110111001001011010101100101001101101110010100000001101; end
            14'd10433 : begin out <= 64'b0010100101000000000111101000111000100101101101000010100001110111; end
            14'd10434 : begin out <= 64'b1010101000000001101010101110000000100010001001011010001110100011; end
            14'd10435 : begin out <= 64'b0010101010111001000111011010101010101001011010011010100001111011; end
            14'd10436 : begin out <= 64'b0001010001110000000110001001001110101010100000011010100010100000; end
            14'd10437 : begin out <= 64'b0010101010011001001010010100010100100010110101100010100101101001; end
            14'd10438 : begin out <= 64'b1010000111001011100111000100101010101001111100101010101001000011; end
            14'd10439 : begin out <= 64'b1010001101101000101010010100001000101011100001011010011110100110; end
            14'd10440 : begin out <= 64'b1010001010000010001001111011101100101001001111111001011000111100; end
            14'd10441 : begin out <= 64'b0010011100100010001010101101010110100111111011100010101001110001; end
            14'd10442 : begin out <= 64'b1010011110101100101010111110110010100111001000111010101010011011; end
            14'd10443 : begin out <= 64'b1010010010000110001010010111100110100101000110001010011110100100; end
            14'd10444 : begin out <= 64'b1010010101001000000111010110010110101011101010111010011001101111; end
            14'd10445 : begin out <= 64'b1001100010011111001000001001010110101010111101100010101011000010; end
            14'd10446 : begin out <= 64'b0010100100011000101001011000101010011100110110001010101101000110; end
            14'd10447 : begin out <= 64'b0010101110011010100101010111101100100100011000100001111011101110; end
            14'd10448 : begin out <= 64'b0010001011001111001010100001110000011000000001001010101010011000; end
            14'd10449 : begin out <= 64'b0010101110011101100111111101100000100101110000010010000010111010; end
            14'd10450 : begin out <= 64'b0010110000001110001010010101011100101010101000001010010111110011; end
            14'd10451 : begin out <= 64'b1001111001001111101010100100011110011101100001100010010001010100; end
            14'd10452 : begin out <= 64'b0010010100010010001000100001001100011001100100110010100000000100; end
            14'd10453 : begin out <= 64'b1010000101101101101010001011100110101010001110010010011000011010; end
            14'd10454 : begin out <= 64'b0010101111010000001010110001110000100001000001101010000011110111; end
            14'd10455 : begin out <= 64'b1010101101001011101010011111011010101010111110110010100101111110; end
            14'd10456 : begin out <= 64'b0010100011110011001001111000110010101000100100101010101111101000; end
            14'd10457 : begin out <= 64'b1010100010000101001010111100101110101001100011001010000011110010; end
            14'd10458 : begin out <= 64'b1010011011111011001001001000010100011101100011111010100111011101; end
            14'd10459 : begin out <= 64'b1010101101011101001010100110101010100100101101110001110111001110; end
            14'd10460 : begin out <= 64'b0010000000011001101010100111010100101000000101100010100110101000; end
            14'd10461 : begin out <= 64'b1010011110110011101010001000001100101001101111000010101101101001; end
            14'd10462 : begin out <= 64'b1010101000100011101001111111001100100100100111111010011111000000; end
            14'd10463 : begin out <= 64'b0010000111110110001001001010011010100100000110101010100000000100; end
            14'd10464 : begin out <= 64'b1001110101001000101010000000101000101100000100110010010010001010; end
            14'd10465 : begin out <= 64'b0010101111110101101001011000110010100110011010000010110000100110; end
            14'd10466 : begin out <= 64'b1010100101100101001001110110011110100010000010111010100110000010; end
            14'd10467 : begin out <= 64'b0010101010100000101010110111101100100101111010011010101100100010; end
            14'd10468 : begin out <= 64'b0010100011011101001001100110001100100110110001110010011001000101; end
            14'd10469 : begin out <= 64'b1010010011110011000110100011000000010000100100010010011111010110; end
            14'd10470 : begin out <= 64'b0010000010000011101010011010010000011111100100000001111110010110; end
            14'd10471 : begin out <= 64'b1001101010100011001001110110111010101000001000101010100101010001; end
            14'd10472 : begin out <= 64'b0001000100011001101001011001110110101000100100101010001001011111; end
            14'd10473 : begin out <= 64'b0010001000110000101010010000100110101001110011111010101010101000; end
            14'd10474 : begin out <= 64'b0010001010111110101010110111010100101001010000000010011011111110; end
            14'd10475 : begin out <= 64'b0010011111000100101010110000100010011010100000111010010000101010; end
            14'd10476 : begin out <= 64'b0010101111010101000111001111001010101011000000011010010111110001; end
            14'd10477 : begin out <= 64'b0010100011010001101010000100101000101000110100110010000110110101; end
            14'd10478 : begin out <= 64'b1001111011001101000110111011000100101010001100101010101111011101; end
            14'd10479 : begin out <= 64'b0010101110000101001010001111101110011011110111111010001101000000; end
            14'd10480 : begin out <= 64'b1010010010001010101010001000110110101011110011110010001000101111; end
            14'd10481 : begin out <= 64'b1010011101000001001000111011101110101000001001101010100110111001; end
            14'd10482 : begin out <= 64'b0001111011110000000110000011101100101011010101001010011101101100; end
            14'd10483 : begin out <= 64'b0000001000011000000111001000101110010011011110001001110001100100; end
            14'd10484 : begin out <= 64'b1010010000110010001001101001101000100111111111111001101111111101; end
            14'd10485 : begin out <= 64'b0010100110111011101010111110011000101010100000000010101000101101; end
            14'd10486 : begin out <= 64'b0001111100001101001001010000000100101011110101000001010001101101; end
            14'd10487 : begin out <= 64'b1010100011011010001010100000101100010010101101101001000111000101; end
            14'd10488 : begin out <= 64'b1001011001101111101000101110110110011000111100101010000100100000; end
            14'd10489 : begin out <= 64'b1010001010000100001010000000000000011101001000001010011011000010; end
            14'd10490 : begin out <= 64'b1010011000010111101010010001111010100111100000111010000110100110; end
            14'd10491 : begin out <= 64'b1010011111101110000111101100001110011110011000011010011111000101; end
            14'd10492 : begin out <= 64'b1010001101000110101010001111100000101011111100101010011011010111; end
            14'd10493 : begin out <= 64'b1010010111011000001000011000001000100000110000111010101000110110; end
            14'd10494 : begin out <= 64'b0010101010110000001001011010111010101010101100011010101111110101; end
            14'd10495 : begin out <= 64'b1010100101011101101010100110011010101010101101010010101111000110; end
            14'd10496 : begin out <= 64'b0001111111011001001010011011101000100100011101011010011011001111; end
            14'd10497 : begin out <= 64'b0010000001100111101001100111100100100100100100111010101000110010; end
            14'd10498 : begin out <= 64'b1010101101010101001010001111010000101010111000101010000101011100; end
            14'd10499 : begin out <= 64'b0010101110000001101010110110011000101010110000110001111100101001; end
            14'd10500 : begin out <= 64'b1010101100010011101010010010101110101000000000000010001011010111; end
            14'd10501 : begin out <= 64'b1010100001110101001001111000111010101010111010010010101000010000; end
            14'd10502 : begin out <= 64'b1010101111010001001010101000110100011011011111111010011110000001; end
            14'd10503 : begin out <= 64'b0010101111111100001001000110011110101001001111000010101111001100; end
            14'd10504 : begin out <= 64'b0010001100110010001000100111110010011101011011001010100100000110; end
            14'd10505 : begin out <= 64'b0010101101100001101010000101111100101010110000110010010001011100; end
            14'd10506 : begin out <= 64'b0010101001001100101010010100110110010001111110101010100000100000; end
            14'd10507 : begin out <= 64'b1010100010011000001001011101011000101010010010110010100001111000; end
            14'd10508 : begin out <= 64'b0010001010010100101001100101101010011111000110001010100000000111; end
            14'd10509 : begin out <= 64'b0010000110101100101010001111101000101010100000100010101011000101; end
            14'd10510 : begin out <= 64'b0010000001101110101001000001100110100001111110101010101001111000; end
            14'd10511 : begin out <= 64'b1010101101100001101010000100100000101010111000101010101110101111; end
            14'd10512 : begin out <= 64'b1001111111101001101000111000100100100100011100111010011100001110; end
            14'd10513 : begin out <= 64'b0010100010001010001001010000011010100101001000001010010000101110; end
            14'd10514 : begin out <= 64'b0010001110010011101010010001101110011110111111011010110000000110; end
            14'd10515 : begin out <= 64'b0010101111001000101001011001110100011101001011100010011010001000; end
            14'd10516 : begin out <= 64'b0010100001111101101010111101110100101010001111110010100001101111; end
            14'd10517 : begin out <= 64'b1010010010010100001010100100110110101001010010101010100000000101; end
            14'd10518 : begin out <= 64'b1010100111100110001001110110111100101011101010011010000111111001; end
            14'd10519 : begin out <= 64'b0010101100100010101010011100110010100111111101111010101100000100; end
            14'd10520 : begin out <= 64'b1010101010101110100101011010000110100101000110100010011110011101; end
            14'd10521 : begin out <= 64'b0010010111100000001010010011110010100111110001111010100110111110; end
            14'd10522 : begin out <= 64'b0010101001111100101001101100101110100110011000100010010000100000; end
            14'd10523 : begin out <= 64'b1010101011011001001010011100101110100001011001110010100010110100; end
            14'd10524 : begin out <= 64'b1010100101111100101001110000101010100011001101011010100000111100; end
            14'd10525 : begin out <= 64'b0010100100011100001001100001101000101010010101010010101010010001; end
            14'd10526 : begin out <= 64'b0010110000111001001010000111011110100100110011101010100101100001; end
            14'd10527 : begin out <= 64'b0010101101010000101010001011111010010101010011111001010110010010; end
            14'd10528 : begin out <= 64'b1010100110110110101010100001000000101000101111000001111110000100; end
            14'd10529 : begin out <= 64'b0010101001101111101010111111101100101010101010001010100110101100; end
            14'd10530 : begin out <= 64'b1001100110101100101010110011111100011011001000101001111001100001; end
            14'd10531 : begin out <= 64'b1010100001001010000111100010000010100001101101100010011100001001; end
            14'd10532 : begin out <= 64'b0010010100100100001010101100011010100011010110111010010110000101; end
            14'd10533 : begin out <= 64'b1010011101100001000101000011010100100110110011001010011011110101; end
            14'd10534 : begin out <= 64'b1010010011001011001010011101000110100110010000000001111110101100; end
            14'd10535 : begin out <= 64'b1010100100011011100111000110010100001011001000011010100111000111; end
            14'd10536 : begin out <= 64'b1010000001000011001000011100001010101010010111010010001010101111; end
            14'd10537 : begin out <= 64'b1010101000100001001000010001010010101010000010101010101000010111; end
            14'd10538 : begin out <= 64'b1010100001101011001011000001011100101000101111000010011000011100; end
            14'd10539 : begin out <= 64'b0010000011011011001010011010000010101010101101001001110110100011; end
            14'd10540 : begin out <= 64'b1010100001101110001000010010001000100010011011011010100111010000; end
            14'd10541 : begin out <= 64'b0010010111001101101010000010001110100110110111010010101100001010; end
            14'd10542 : begin out <= 64'b1010011001011000101010100100011100101010010101111010011010010110; end
            14'd10543 : begin out <= 64'b1010011001100011001010100110001010101000010010101010101011010001; end
            14'd10544 : begin out <= 64'b1010100000111011100111110001001010100100110011000010010111011000; end
            14'd10545 : begin out <= 64'b1010000110001111101001111110011000100010011110001010100011011111; end
            14'd10546 : begin out <= 64'b1010110000000011101001001010100100100100101111100010100111010011; end
            14'd10547 : begin out <= 64'b1010100010101011101001111010110100101000100010010010000000001011; end
            14'd10548 : begin out <= 64'b1010011110101100001001010100011110101010101000011010000111011100; end
            14'd10549 : begin out <= 64'b1001100101101011001001100110101010100000011101011010101101110000; end
            14'd10550 : begin out <= 64'b0010000101010111101001011011101000101011111101001010001011000000; end
            14'd10551 : begin out <= 64'b1010101010101000101010010000001010101001101001001010000011010100; end
            14'd10552 : begin out <= 64'b1010101110001110001000111010110010101001111100100010101001111110; end
            14'd10553 : begin out <= 64'b1010010100101100001001111101010100100111000110001010010000100010; end
            14'd10554 : begin out <= 64'b1010100101011100001010110000000010101010111100111010011010011110; end
            14'd10555 : begin out <= 64'b1010100001101001101001101010010010100101110011001010101100101101; end
            14'd10556 : begin out <= 64'b0010010101001010001010110101001000101001100100101010100110101000; end
            14'd10557 : begin out <= 64'b1010100101100111101010000111101010101010111111100010001000001001; end
            14'd10558 : begin out <= 64'b1010101110001011001001101100001010100100001001110010100010011010; end
            14'd10559 : begin out <= 64'b1010001001101110001010010001101100101010110110001010101100001010; end
            14'd10560 : begin out <= 64'b0010100110000010101010111101001010101011100111101010010111000001; end
            14'd10561 : begin out <= 64'b0010100001011001101001001001101100101010000101010001111111001000; end
            14'd10562 : begin out <= 64'b1010010101011011001010100110000100100001101100000010010110101110; end
            14'd10563 : begin out <= 64'b1010010101001000001010110001010110101010100100000010011011111001; end
            14'd10564 : begin out <= 64'b0010010101010100001001000110111100101000100001100010100111010100; end
            14'd10565 : begin out <= 64'b0010001010101010001010010110011100100000100010101010010110100101; end
            14'd10566 : begin out <= 64'b1010100110111011001010000001110100101011010100100010100101001001; end
            14'd10567 : begin out <= 64'b0010001101010010001010001100101010100000001101000010100110001101; end
            14'd10568 : begin out <= 64'b0010011100000111001010000111011000101001101001001010010011001000; end
            14'd10569 : begin out <= 64'b1010101011000111001010110001001100101000010010010010010100111111; end
            14'd10570 : begin out <= 64'b1001111011001010101010111111000000011000001010001010000101001011; end
            14'd10571 : begin out <= 64'b0010010001100100001001101010111000100000100110101010000100011111; end
            14'd10572 : begin out <= 64'b1010010001000100100100111010011010100111111110001010010011100010; end
            14'd10573 : begin out <= 64'b1010011001011000101010110111010100101001000100111010100010101101; end
            14'd10574 : begin out <= 64'b1010101110101010001010011110000110101001001011111010001111101000; end
            14'd10575 : begin out <= 64'b1010100000011111001010110110011110011101110110000010101110011101; end
            14'd10576 : begin out <= 64'b0010010111100010000111100011111100101001010101110010100111001010; end
            14'd10577 : begin out <= 64'b0010000001000001001000100011111000101010011010110010010010000100; end
            14'd10578 : begin out <= 64'b1000110000100110001001010001100000100011101000001010100000100001; end
            14'd10579 : begin out <= 64'b0010010011100110001011000000100010101000111101101010010001101111; end
            14'd10580 : begin out <= 64'b1010010110001001001010111100011000101011101111010010101001000111; end
            14'd10581 : begin out <= 64'b1010010111100010101010110000000100100111100010001010100001100110; end
            14'd10582 : begin out <= 64'b0010010100111010000111111010001100100101010111010010011010100111; end
            14'd10583 : begin out <= 64'b0010010111110110101010001111111110101011111000111010101111010101; end
            14'd10584 : begin out <= 64'b1010100001111110001010010011100100101010010100001010101110010000; end
            14'd10585 : begin out <= 64'b1010101100010010101001100000010010101001000000101001010000010001; end
            14'd10586 : begin out <= 64'b0010101001001001101010110101111100100001110101000010011001010000; end
            14'd10587 : begin out <= 64'b0010010001011000001000001100001100100011010000100010011010111010; end
            14'd10588 : begin out <= 64'b0010101111001101101000110101010000100111000001001010100101100001; end
            14'd10589 : begin out <= 64'b1010011111101010001010010000011010101011111111010010001011001001; end
            14'd10590 : begin out <= 64'b0010100101110100101010001000101110101010100111100010101110010110; end
            14'd10591 : begin out <= 64'b0010100011110110001000100111100110100111111010110010101101011111; end
            14'd10592 : begin out <= 64'b1010100110111001101000011111010000100001000000001010100101110110; end
            14'd10593 : begin out <= 64'b1001111010011110101001110011011010100101011110001010011010101010; end
            14'd10594 : begin out <= 64'b0010011100111011001000110111101000011011000111110010101010100011; end
            14'd10595 : begin out <= 64'b1010101010111100001001110011101110101000011101101010000100111001; end
            14'd10596 : begin out <= 64'b0010101011100101101010110110001000101010010000101010101100101100; end
            14'd10597 : begin out <= 64'b0010101110101011000111001100011110100010110011101001111101101101; end
            14'd10598 : begin out <= 64'b0001111100011001001010011000000100100110010100000010101110000110; end
            14'd10599 : begin out <= 64'b1010011100000001101001011111100000101001011000010010100110111101; end
            14'd10600 : begin out <= 64'b0010100101100011001001100111100010101001000010001010011001011011; end
            14'd10601 : begin out <= 64'b1010101001001001101010010110010110100110010110000001110011011111; end
            14'd10602 : begin out <= 64'b0010101111010110101001011110010100101010001110101010001011011100; end
            14'd10603 : begin out <= 64'b0010000101011010001010000011111010101001000000000010001101110101; end
            14'd10604 : begin out <= 64'b0010100000000110001001101111010000101001101101010010100101000100; end
            14'd10605 : begin out <= 64'b1001100010010111001010010110101110011000010101111010001110001000; end
            14'd10606 : begin out <= 64'b1010011011101111001001000010000010010111011110110010101001011000; end
            14'd10607 : begin out <= 64'b1010000100001010000101001000010110100000111000010010100010010010; end
            14'd10608 : begin out <= 64'b0010100011110011101010010000110110101000010010001010001001000000; end
            14'd10609 : begin out <= 64'b1010100111110110001010000110000010100010001000000010100010010000; end
            14'd10610 : begin out <= 64'b0010100001111010101010110000011110100100001001010010100000110110; end
            14'd10611 : begin out <= 64'b1010011100101101101010110011010100101000101010010010101010110000; end
            14'd10612 : begin out <= 64'b0010001101001011001001110101000000101000101000011010010101000111; end
            14'd10613 : begin out <= 64'b0010101001011010101001010011100010011110001001100010100000010110; end
            14'd10614 : begin out <= 64'b0010010111010111101000011111011010001110010111111010010010000100; end
            14'd10615 : begin out <= 64'b1010101001001101101000000011000110101011011111010010001101010111; end
            14'd10616 : begin out <= 64'b0010101011100011001010110011110000101001100101101010000011111011; end
            14'd10617 : begin out <= 64'b1010100000011111001001101100100010100001000110100010100110111000; end
            14'd10618 : begin out <= 64'b1010010011000100000110101010100100101011000110010001111101101111; end
            14'd10619 : begin out <= 64'b1001111000001010101000111111011010101001010000000010110000001100; end
            14'd10620 : begin out <= 64'b0010001110011010101010001000011110100110010001101010101111101001; end
            14'd10621 : begin out <= 64'b0010100100011110101010100100111000100110000110000010101101101011; end
            14'd10622 : begin out <= 64'b1010011110001100001000101010111010100101111011001010101111001011; end
            14'd10623 : begin out <= 64'b1010100110011100101010011010010100100100001100100010001110001111; end
            14'd10624 : begin out <= 64'b1010011000100011001001101101111000101010101001110010100111110111; end
            14'd10625 : begin out <= 64'b0010010000101111101001001011000110100110110001110010110001100001; end
            14'd10626 : begin out <= 64'b1010101100101011101001110110110000100101010111100010000010101111; end
            14'd10627 : begin out <= 64'b1010001010110010000110001110101110101000101000111001110111011001; end
            14'd10628 : begin out <= 64'b1001111111001011001001001111100100101001111010111010101010101110; end
            14'd10629 : begin out <= 64'b1010101000001011101000010001110100101010011000101010101100000101; end
            14'd10630 : begin out <= 64'b0010010101110101101001110011100010100001110101011010000110010111; end
            14'd10631 : begin out <= 64'b0010101111101100101010110000010000100101110111110010100100001010; end
            14'd10632 : begin out <= 64'b1010100001110110101010100100111000101011101001100001100010001100; end
            14'd10633 : begin out <= 64'b0010100111010110100100011100000010100100100001111010100111111000; end
            14'd10634 : begin out <= 64'b0001100101100011000110110011001010100001110001111010100010011001; end
            14'd10635 : begin out <= 64'b1000111011000111001000010000110100101010110010111010101111001001; end
            14'd10636 : begin out <= 64'b0010011111111100001001101101000100100100001110101010101001001011; end
            14'd10637 : begin out <= 64'b1010101101011110101010110100101010100010000101011010101110011010; end
            14'd10638 : begin out <= 64'b1010100001100110001010111100010110011001111100101010100010010000; end
            14'd10639 : begin out <= 64'b1010100110010000001010110100000100101000001001101010101110001000; end
            14'd10640 : begin out <= 64'b0010010000110011001001111111001000101000001010010010011010010001; end
            14'd10641 : begin out <= 64'b0000000000100011001001000000100100100101011110100010101100101011; end
            14'd10642 : begin out <= 64'b1010101011110111001000001000001010101011111011100010000110100010; end
            14'd10643 : begin out <= 64'b1010100101011000101001101101010110100001001010011000100101110100; end
            14'd10644 : begin out <= 64'b0010010001111011101010100001100110100000001100110010001101110100; end
            14'd10645 : begin out <= 64'b0010101001011001001001010010101000100101010011000010101010100000; end
            14'd10646 : begin out <= 64'b1010101010011100001010010010101100101001111111111001111100001000; end
            14'd10647 : begin out <= 64'b0001111010111001001010010011001000100100111000000010100011011000; end
            14'd10648 : begin out <= 64'b1010100011100100001001100001100010101001011110010010010101111001; end
            14'd10649 : begin out <= 64'b1010101001010110100110110111100010101000111010000010001110000110; end
            14'd10650 : begin out <= 64'b0010100111101110100101010010001000011101110011011010011100010001; end
            14'd10651 : begin out <= 64'b1010011001100110101000011010010110101000010110001010100101011000; end
            14'd10652 : begin out <= 64'b0010100100000101101010110001100010100000100100000010010101111100; end
            14'd10653 : begin out <= 64'b1010101111000001000110111001010110100010101101000010101100110000; end
            14'd10654 : begin out <= 64'b0001101100110110001010011011111100100101011110100010100010011101; end
            14'd10655 : begin out <= 64'b0001110000010111101001010010110010100011101000101010101110110101; end
            14'd10656 : begin out <= 64'b1010101011000001101010001111001110100100011001000010011011011000; end
            14'd10657 : begin out <= 64'b0010100100110101001010100100001100100000100101110010100111000000; end
            14'd10658 : begin out <= 64'b0010100001011010001010001011100000101001010011111010110000001110; end
            14'd10659 : begin out <= 64'b1010011110000100101010001100000000101010100100010010011101101100; end
            14'd10660 : begin out <= 64'b1010101011100011101001111101110100011010111001011010100110000100; end
            14'd10661 : begin out <= 64'b0010100011110100001001010101010100101001001110011010010000111000; end
            14'd10662 : begin out <= 64'b1010100101010011100111000101101110100111100000000010100011010010; end
            14'd10663 : begin out <= 64'b1010011110001010001000011010100010100010010011010010101111101110; end
            14'd10664 : begin out <= 64'b1010101010111001001010100001010000011101010010110010101011101000; end
            14'd10665 : begin out <= 64'b0010100011100011001010000010110010100100100011001010100101100100; end
            14'd10666 : begin out <= 64'b1010011001001100101001100010011100100100001110110010000010101011; end
            14'd10667 : begin out <= 64'b0001010100111100001001101000110100100000111100101010011001000001; end
            14'd10668 : begin out <= 64'b1010110000001100101010001111101110100011011011101010100101010110; end
            14'd10669 : begin out <= 64'b1010100010011000001001111010001110100110010010110001110111100100; end
            14'd10670 : begin out <= 64'b1010000110011000001010100110001110010111101001011010101000010011; end
            14'd10671 : begin out <= 64'b1010001101101010101010111110111110011110010000110001111000010010; end
            14'd10672 : begin out <= 64'b1010001011110100001001110010101110101000001011000010100100100001; end
            14'd10673 : begin out <= 64'b1010000101000010001001110011010010101000011010001010001010001011; end
            14'd10674 : begin out <= 64'b0010101011101101000111111100100000100100100111011010101100000111; end
            14'd10675 : begin out <= 64'b1010100100010011101001111010100000101000011001101010011101001000; end
            14'd10676 : begin out <= 64'b1010101110111110001010111001000110100100100001101010101110000010; end
            14'd10677 : begin out <= 64'b1010010101100110101000110011001100011000111101111010000001000010; end
            14'd10678 : begin out <= 64'b1010010100111011101010101001111000010111001101100010010000110100; end
            14'd10679 : begin out <= 64'b1010101101010000001010000101010110101011011110101010011011010100; end
            14'd10680 : begin out <= 64'b1010100110000011101010110101010100011110101100100010100011100110; end
            14'd10681 : begin out <= 64'b1010000100111000001000010110100100100000001101111010100111100010; end
            14'd10682 : begin out <= 64'b0010100010010000001010000001111110101011011101011010010011001100; end
            14'd10683 : begin out <= 64'b0010101101011001101010101010110010101001101111001001011011000011; end
            14'd10684 : begin out <= 64'b0010010001000100100110100101010110011101111010010010010000110110; end
            14'd10685 : begin out <= 64'b1010011100100010101010001111000100101001100110111010100001100010; end
            14'd10686 : begin out <= 64'b1010100011000011001001111100101010100100010010001010101101000011; end
            14'd10687 : begin out <= 64'b0010100010001101100111001110101100101010100011011001110011101000; end
            14'd10688 : begin out <= 64'b0010100011101001001010110000000100101010100100100010011000101010; end
            14'd10689 : begin out <= 64'b0010101000010000101000111111111010100100001001100010101100111001; end
            14'd10690 : begin out <= 64'b1010101001110111001010001110011110100000000011010010100010100110; end
            14'd10691 : begin out <= 64'b0001110100011101101010000100110000101010110001111010100000000110; end
            14'd10692 : begin out <= 64'b1010000000100111101010101010100110100110010111000010010110111110; end
            14'd10693 : begin out <= 64'b0010101011010010101011000001010000101000111000100010000101010000; end
            14'd10694 : begin out <= 64'b0001111111010110101010001010010010101001000010110010100001101001; end
            14'd10695 : begin out <= 64'b1001110011100101101010001011000010101000000010011010101010111001; end
            14'd10696 : begin out <= 64'b1001111100010000001001110100110110011111111011111010100011101000; end
            14'd10697 : begin out <= 64'b0001101110100110000101111111101000101010111110000010011010010000; end
            14'd10698 : begin out <= 64'b0010011110001011001000111111001010101010110001000010101001010000; end
            14'd10699 : begin out <= 64'b1001100010010111101010001001011010011110101011100010010000000010; end
            14'd10700 : begin out <= 64'b0010001000111111101001011000000110011001111111110001110111111101; end
            14'd10701 : begin out <= 64'b1010010010010100001001011010110000100100011001110010011101111010; end
            14'd10702 : begin out <= 64'b1001101101101000101000100110011010101010001100011010100111101101; end
            14'd10703 : begin out <= 64'b0010101101101100001010111111111010101000110011111010100111000011; end
            14'd10704 : begin out <= 64'b0010101111111001101010100110110010101000001101101010101100001010; end
            14'd10705 : begin out <= 64'b1001110010001011101000111110110110101000010010000010110000001101; end
            14'd10706 : begin out <= 64'b0010000110110100001000011001111010100011100011000010110001101110; end
            14'd10707 : begin out <= 64'b1010101111011011101010101001000100100100100101001010101110100000; end
            14'd10708 : begin out <= 64'b1010101101111110101001011101101010100101011000111010010101011001; end
            14'd10709 : begin out <= 64'b1010100011100001001000100011101010010001000110101001101001101111; end
            14'd10710 : begin out <= 64'b0010001110110110001010010101110000101011100101001010100111010001; end
            14'd10711 : begin out <= 64'b0010100111000001001001111000100110100101000001110010100001100001; end
            14'd10712 : begin out <= 64'b1010100111011001001010100011101010101001010111110010010101010101; end
            14'd10713 : begin out <= 64'b0010010000001100101010000011101110100110111110100010001001101000; end
            14'd10714 : begin out <= 64'b1010010010010100101010100000000000100110001001011010100101100010; end
            14'd10715 : begin out <= 64'b1010010001010010001001001100011110011011000100010010100100101100; end
            14'd10716 : begin out <= 64'b0010100100101111101001000000110100010101110101101010010011101100; end
            14'd10717 : begin out <= 64'b0010011000100110100111001110111100100100010010111010001111011100; end
            14'd10718 : begin out <= 64'b0010100111001000101010010100110100101001110010011010101011100101; end
            14'd10719 : begin out <= 64'b0010010000100100001010100001010010101010001101101010101000100010; end
            14'd10720 : begin out <= 64'b1010010100101100101010010100011000100000110111111010011011000011; end
            14'd10721 : begin out <= 64'b1010100100011110001010110101000010100110011001000001111111110010; end
            14'd10722 : begin out <= 64'b0010010001100001101010100100101110101010110110101010101000110010; end
            14'd10723 : begin out <= 64'b1010101011101001101001000100110100101001101001011010010111000001; end
            14'd10724 : begin out <= 64'b0010100101101111101010000110110010101011000011001010101111011001; end
            14'd10725 : begin out <= 64'b0010101010110100101010110001100100101010010101101010011000111111; end
            14'd10726 : begin out <= 64'b0010100111111010101000111011110000101001110010011010101000011011; end
            14'd10727 : begin out <= 64'b1010010111111111001000001101001000101000011000111010101011100100; end
            14'd10728 : begin out <= 64'b0010100011000111001010011100101000101010100000111010101011010011; end
            14'd10729 : begin out <= 64'b0010010001111000001010100111110000100000101001011010101001000110; end
            14'd10730 : begin out <= 64'b1010100100011110100111111111000100001011001001110010101000110001; end
            14'd10731 : begin out <= 64'b0010001111101000001010010001001000100100010101100010001101101010; end
            14'd10732 : begin out <= 64'b0010100110000100001010001101111000101010111010100010100111000000; end
            14'd10733 : begin out <= 64'b1010010011100100001010100100101100101001111111101010101000101111; end
            14'd10734 : begin out <= 64'b0010100110111001001010110110100110101011000011010010100000011110; end
            14'd10735 : begin out <= 64'b1010101110001101001001101101011110011000010011000010101101000101; end
            14'd10736 : begin out <= 64'b1010100111001000101000011011100000011010010010000010101100110101; end
            14'd10737 : begin out <= 64'b0010101101000010101010111111011000100111100111000010100111001011; end
            14'd10738 : begin out <= 64'b0010001010010110001010011011011010101000110101010010010010111010; end
            14'd10739 : begin out <= 64'b1010100101111110101000111100000100100011010001100010100000010001; end
            14'd10740 : begin out <= 64'b0010101100010001001010010110001110101000100110000010101101001011; end
            14'd10741 : begin out <= 64'b1010000111100100001001101110001000011010110111100010011010000011; end
            14'd10742 : begin out <= 64'b1010011101001010101001001001001100101001010111010010100100000000; end
            14'd10743 : begin out <= 64'b0010011000000000001001110111011100011110110110011001101011101010; end
            14'd10744 : begin out <= 64'b1010101000001101101001101010010100010010010100010010100111110101; end
            14'd10745 : begin out <= 64'b1010100110100001000111011000010010011111100000100010100111001100; end
            14'd10746 : begin out <= 64'b0010100011110100101010010111010110011001000101100010100111001010; end
            14'd10747 : begin out <= 64'b0010100001110000001010110101001100101010011010010010100001001001; end
            14'd10748 : begin out <= 64'b0010100111101000101001000111000110101000111101010010100101111110; end
            14'd10749 : begin out <= 64'b1010011001110010101001001111100000101010011110001010011101110110; end
            14'd10750 : begin out <= 64'b0010010100111101001011000000011000101011110010110010101111111001; end
            14'd10751 : begin out <= 64'b0010011101100110101001011100000100101001100100000010101011000011; end
            14'd10752 : begin out <= 64'b0010101000111010001001100101110010100000000010100010100000100000; end
            14'd10753 : begin out <= 64'b0010010100001000101001001111011000101000101110011010100100101110; end
            14'd10754 : begin out <= 64'b1001111011111101001010110000001000101001011000111010101111001011; end
            14'd10755 : begin out <= 64'b1001010000110011101010010011001000011001000011110010000101110010; end
            14'd10756 : begin out <= 64'b1010101001010010101010011001111100101010101101001010100110001111; end
            14'd10757 : begin out <= 64'b1010101011011010100110001000010110010011100000110010100010011001; end
            14'd10758 : begin out <= 64'b0010100100000101000111000000010010100111110001011010010010101110; end
            14'd10759 : begin out <= 64'b0010110000010101001001101011010110100101100100001010100001010001; end
            14'd10760 : begin out <= 64'b1001110011010011101010110111000000100010001110111010000000010111; end
            14'd10761 : begin out <= 64'b0010010110101000101010110100101100100011110011001010101010101000; end
            14'd10762 : begin out <= 64'b0001111011010101000110000011000100101010110000101010100111000000; end
            14'd10763 : begin out <= 64'b0010100010110000001010101100011000011111110000101010011010110000; end
            14'd10764 : begin out <= 64'b0010000010111000001010101110001010101001011111010010100000011001; end
            14'd10765 : begin out <= 64'b0010101111000111101001100010110100100110010101110010101001001101; end
            14'd10766 : begin out <= 64'b0010100001101001001010001010011110101010010111101010100101101111; end
            14'd10767 : begin out <= 64'b0010010100010001101010011010010000101010100100000001110101000010; end
            14'd10768 : begin out <= 64'b0001111111101010101001111000100000101000101110100010101111110110; end
            14'd10769 : begin out <= 64'b1010101000010011101001010001011110100001110110110010100011010101; end
            14'd10770 : begin out <= 64'b0010011011011010001001111101010010101010110101110010000100011011; end
            14'd10771 : begin out <= 64'b1001110001001010000111000000001110101000111111110001010001111000; end
            14'd10772 : begin out <= 64'b0010100011011000101010010011110100101001101101010010101010111111; end
            14'd10773 : begin out <= 64'b1010000011011110101001011100100100100011000110010010101000110010; end
            14'd10774 : begin out <= 64'b1001111001001110101001100100100110100010000100101010101110100110; end
            14'd10775 : begin out <= 64'b1010001100011011001010111101111100100010001111001010011110010010; end
            14'd10776 : begin out <= 64'b1010000110010100101000111101110110101010100111011010001111100110; end
            14'd10777 : begin out <= 64'b0010101101011110101001110100111010101011010000010010010011111000; end
            14'd10778 : begin out <= 64'b1010010101111111001010010101111100101001000010000010100011110010; end
            14'd10779 : begin out <= 64'b1010100110100000101010101100111100101000101000010010010111010101; end
            14'd10780 : begin out <= 64'b0001110110110100101010100111000100101010011101110010011000000010; end
            14'd10781 : begin out <= 64'b0010100011100100000111100001110000101000111010011010100010110101; end
            14'd10782 : begin out <= 64'b0010100100001011001001110111000010101000010111001010101011010111; end
            14'd10783 : begin out <= 64'b1010011101000010101001100010101110100110001001000010100111101010; end
            14'd10784 : begin out <= 64'b0010011000110010001010001010100010101010011101011010100100101110; end
            14'd10785 : begin out <= 64'b0001111111101111000111111100000010100111000100101010100001100111; end
            14'd10786 : begin out <= 64'b1010100000001110001010011000100110101010110010101010101000101110; end
            14'd10787 : begin out <= 64'b1010001010011001101001101101000100101011010101000010100100000110; end
            14'd10788 : begin out <= 64'b1010011110010011001010100111011000101010111010110010100110100011; end
            14'd10789 : begin out <= 64'b0010101001111101001010111110101000100101100011111001100110001111; end
            14'd10790 : begin out <= 64'b0010011111010110001010011000110100101010101101110010100011001011; end
            14'd10791 : begin out <= 64'b1010100100011010100111010101010000100111110100011001101110111001; end
            14'd10792 : begin out <= 64'b1010101001010000001001001001100000101010111110001010101010110111; end
            14'd10793 : begin out <= 64'b1010101100101010001010001011000100100010011101010010100001010100; end
            14'd10794 : begin out <= 64'b1010100101010110001010001111110010011000110101101010010101011110; end
            14'd10795 : begin out <= 64'b0010100001010101001001000010010010100111100100001001011101001011; end
            14'd10796 : begin out <= 64'b1010011101010001001000011011100010011100011000100010010000010000; end
            14'd10797 : begin out <= 64'b1010100101010010100111110010010100101011000101011010100100000011; end
            14'd10798 : begin out <= 64'b1010011111001110101010101111010000100111111100010010011110111001; end
            14'd10799 : begin out <= 64'b1010101001101101101010111110000010101001100000100010101000001100; end
            14'd10800 : begin out <= 64'b0010101011011111001010101100100110010110110000111010101011010110; end
            14'd10801 : begin out <= 64'b0010010000101111100010001110010000101000110110010010010111111110; end
            14'd10802 : begin out <= 64'b0010011110101111001001001100001010011000010100100010010010101011; end
            14'd10803 : begin out <= 64'b1010000100101111001001011000000100100111111010110010100111100011; end
            14'd10804 : begin out <= 64'b1010100101010100101000111010100010101011100010001010100110111101; end
            14'd10805 : begin out <= 64'b1010100101100101001010001111101010100100010010010001001010001100; end
            14'd10806 : begin out <= 64'b0010100110111100100111111011100100011100100000010010101110100100; end
            14'd10807 : begin out <= 64'b0010100011101110101010010110000110101010001001000010101010011111; end
            14'd10808 : begin out <= 64'b1010001010111011101010101000000100100100101000000010010110101110; end
            14'd10809 : begin out <= 64'b0010101000000100101010110101110010101010110011100010011011100000; end
            14'd10810 : begin out <= 64'b0010100100100000101010110001100100101001100101011010011011010000; end
            14'd10811 : begin out <= 64'b1010000000110011101010000100000100100101111001000010100110011001; end
            14'd10812 : begin out <= 64'b0010000101101100100100010110101010101001010001110010101110000000; end
            14'd10813 : begin out <= 64'b0010010110011101101010111101001100100111111000000010011111011111; end
            14'd10814 : begin out <= 64'b0010100001100110001001111010101110101001111000100010101011100010; end
            14'd10815 : begin out <= 64'b0010100011001010001001011011001010101010111011010010100001101010; end
            14'd10816 : begin out <= 64'b1010000100010111001001111111000110101000100000011010100001011111; end
            14'd10817 : begin out <= 64'b0010101011011111101010001110110110101000101011101010011101001010; end
            14'd10818 : begin out <= 64'b1010100111101001101001010110000010101010110100100001111100100000; end
            14'd10819 : begin out <= 64'b1010100010101101000111000111100010100111110011111010101001111110; end
            14'd10820 : begin out <= 64'b1010100001100010100101101011110100101000101100111010001011111110; end
            14'd10821 : begin out <= 64'b0010010100010100101010100001111000101010001000111010100111101100; end
            14'd10822 : begin out <= 64'b1010001011011011101010001110011000101000111000010010011110111100; end
            14'd10823 : begin out <= 64'b1010101111011001001001011010111110101000100110110010010110001000; end
            14'd10824 : begin out <= 64'b1010101101100100101000110110100000101011111011001010011111000110; end
            14'd10825 : begin out <= 64'b1010000100101111101010100011110100100111000011111010101011011110; end
            14'd10826 : begin out <= 64'b1001110000010010101001101000101110101000010011000010010000100010; end
            14'd10827 : begin out <= 64'b1010011001100000001010010011100000010011110100111010011010111100; end
            14'd10828 : begin out <= 64'b0010100101000110101001110100111110101011100001100001111000100101; end
            14'd10829 : begin out <= 64'b1010101101000100100110011100110100101011000101000010011100010111; end
            14'd10830 : begin out <= 64'b1010101111110100101001110001101000100011100000100010100011100000; end
            14'd10831 : begin out <= 64'b1010100011010111101010000000010110010000011101011010011010011101; end
            14'd10832 : begin out <= 64'b0010100011001010101010101100000000101000000111001010101100100101; end
            14'd10833 : begin out <= 64'b1010011000001000000110111101011110011111000010110010100101001100; end
            14'd10834 : begin out <= 64'b1010100010001001100110010111001100101010010001011010000011000100; end
            14'd10835 : begin out <= 64'b0010011110011110101010000100001010101011100011101001110110001101; end
            14'd10836 : begin out <= 64'b1010101001010111001010000101111010101010101010100010000000110001; end
            14'd10837 : begin out <= 64'b1010011000110100001000001100001000101010001100011010001100101100; end
            14'd10838 : begin out <= 64'b1010100101010010001010000000110110100100111100010010100110000000; end
            14'd10839 : begin out <= 64'b0010011100011101001001101101101000101000010101110010100010010000; end
            14'd10840 : begin out <= 64'b0010100111010111001010000111111100101001011011110010101111001110; end
            14'd10841 : begin out <= 64'b0010010110011101001001011101001100100100000011010010100110111001; end
            14'd10842 : begin out <= 64'b1010100000100110101010000000101010101011000000110010011101100001; end
            14'd10843 : begin out <= 64'b1010100110000000100111001001010100101010110110101010100110110011; end
            14'd10844 : begin out <= 64'b1010100000000010100101001010011000101011001111001010011010100111; end
            14'd10845 : begin out <= 64'b1010101000001011101010010100011000011000100111000010100011010010; end
            14'd10846 : begin out <= 64'b1010100010011100001001001110101110100100111111001010010111100101; end
            14'd10847 : begin out <= 64'b1010010010001000101001111101010110100111101010010010010010000111; end
            14'd10848 : begin out <= 64'b1010101110011001001001101011100000101001011101111010100101100101; end
            14'd10849 : begin out <= 64'b0010010010001001001010000001100110100101111001101010011100101001; end
            14'd10850 : begin out <= 64'b0010011000010010001000000110111110100111101111111010010101111111; end
            14'd10851 : begin out <= 64'b0010011100011101101001111100011000101000110111001001100001110100; end
            14'd10852 : begin out <= 64'b1010101001111101101010101001111000101000011011101010010010011110; end
            14'd10853 : begin out <= 64'b0010101111111011001010101001101010101010001110001010011000001110; end
            14'd10854 : begin out <= 64'b1010110000000011101000111100101110011110111110000010100100110100; end
            14'd10855 : begin out <= 64'b1010000111111010100111000000111010101011010010011010010101110010; end
            14'd10856 : begin out <= 64'b1010100011010110100111001001001010101010011110111010100100011010; end
            14'd10857 : begin out <= 64'b0010010101000101101010000110010100101000011101001010010100100110; end
            14'd10858 : begin out <= 64'b0010011010110001001010011101111010101011100110011010101101110101; end
            14'd10859 : begin out <= 64'b1010010100000101101010111000000010100001110100001010100101001010; end
            14'd10860 : begin out <= 64'b1010101111111110101010111010001110101010001101001001100000111101; end
            14'd10861 : begin out <= 64'b0010101100101001001001100011001100100101000000001010100011111001; end
            14'd10862 : begin out <= 64'b0010010010111011101010100000100010101011111010000010011000000101; end
            14'd10863 : begin out <= 64'b0010100010001000001010101001001100100010000000001010101000011010; end
            14'd10864 : begin out <= 64'b1010100010010011001001100001100010010110000001100010100010001111; end
            14'd10865 : begin out <= 64'b0001111101010000100110100101111100011001010110000010010000100010; end
            14'd10866 : begin out <= 64'b0010000101001100100111001001101110100111001110011001111010101000; end
            14'd10867 : begin out <= 64'b0010101001001100100110100010100000101011010000111010011100000100; end
            14'd10868 : begin out <= 64'b0010000010011110001010101111011010100111100010101010010101101101; end
            14'd10869 : begin out <= 64'b0010101001000000001000101111100010011011001101011010100101100010; end
            14'd10870 : begin out <= 64'b1010011010101011001001010110010110011010110100000010100100000010; end
            14'd10871 : begin out <= 64'b0010101000100110101001000110000100101001000011100010011000100111; end
            14'd10872 : begin out <= 64'b0010000101011010001010111011110000101010011100000010000111100011; end
            14'd10873 : begin out <= 64'b1010100011011000001010110000000000101000000000100010011110110001; end
            14'd10874 : begin out <= 64'b0010001010001011001010001111111000100111111001101010101001110110; end
            14'd10875 : begin out <= 64'b0010101000011011101000000000000100101011100101110010100011010000; end
            14'd10876 : begin out <= 64'b0010000000000111001010101101011100100110110110101010100010000101; end
            14'd10877 : begin out <= 64'b0001110000010100001010100000010100101011011000100010011000011111; end
            14'd10878 : begin out <= 64'b0010100010010001101010011011111100100010111000111010010110010011; end
            14'd10879 : begin out <= 64'b0010001001101111100101011010001010001100101101010010100110010001; end
            14'd10880 : begin out <= 64'b0010100010110111001010101010110100100111111101000010101110000000; end
            14'd10881 : begin out <= 64'b0010001000001101001010100101100000100100101011010010101011101011; end
            14'd10882 : begin out <= 64'b1010100011001001001010101110100010100001111011101010010101010001; end
            14'd10883 : begin out <= 64'b1010101011011001001001010000001010010101010010101010001110011100; end
            14'd10884 : begin out <= 64'b0010100000110101101001000001101110101001100110000010101100010110; end
            14'd10885 : begin out <= 64'b1010101000100000101010101011000000101011000000110010101000100101; end
            14'd10886 : begin out <= 64'b1010101100110000101010101111111100101100000011010010011110110011; end
            14'd10887 : begin out <= 64'b1010011010111001001010010101111000011110001010111010101110100000; end
            14'd10888 : begin out <= 64'b1001010010010010101001111000010100010100100001010010100000011100; end
            14'd10889 : begin out <= 64'b1010000010011101001001001101011010011101101001011010011010100010; end
            14'd10890 : begin out <= 64'b1010101001100100001010011001100000101000010101010010011110101111; end
            14'd10891 : begin out <= 64'b1010011000000011001001111001010000100100011111101010001111011010; end
            14'd10892 : begin out <= 64'b1010010111010000001010110001111100100100100010111010011011100010; end
            14'd10893 : begin out <= 64'b1010010111110010001000101101111110101011100101001010001101101100; end
            14'd10894 : begin out <= 64'b1010100111011110101000100000110010100101101011011010101101001010; end
            14'd10895 : begin out <= 64'b1010000110010110101001101100001010101000010111110010101111001110; end
            14'd10896 : begin out <= 64'b1010010000001101001001000000111010101001000001011010001101111101; end
            14'd10897 : begin out <= 64'b1010001100111100101010101010010100101000100110011010101000111100; end
            14'd10898 : begin out <= 64'b0010101001111000101010100000010010101010010100010010100101111101; end
            14'd10899 : begin out <= 64'b1010011100110100100111110111000000101000011100110010100000101101; end
            14'd10900 : begin out <= 64'b0010101110011101101010000011001110101001010011111010101100011101; end
            14'd10901 : begin out <= 64'b0001111000011110001010101011111010100111011101010010100001011111; end
            14'd10902 : begin out <= 64'b0010100100111010001000001100001110101000000001111001110000001111; end
            14'd10903 : begin out <= 64'b1010010111011011101010011010001010100110011111000010100011010101; end
            14'd10904 : begin out <= 64'b0010100010011110101000111101101110100111100111001010100000100100; end
            14'd10905 : begin out <= 64'b1010010111000111001001011000101110100010111001110010100011011001; end
            14'd10906 : begin out <= 64'b1010001011100111001010101011101000100011101101000010100101010111; end
            14'd10907 : begin out <= 64'b1010110000000001101000100010110100101001111111010010101100010110; end
            14'd10908 : begin out <= 64'b1010101010011111101001011000110110100111101110001010011100001111; end
            14'd10909 : begin out <= 64'b1010100000101100101010011011100100101010110110100010011010110001; end
            14'd10910 : begin out <= 64'b0010101000001001001000011110101100100100110010010010001000000101; end
            14'd10911 : begin out <= 64'b1010001101011010001010110001000000101000011111001010001100101101; end
            14'd10912 : begin out <= 64'b0010011111010111000111111101000010011110010011010010010111000111; end
            14'd10913 : begin out <= 64'b0001110111100001001010001101011110101011101110000010101100001100; end
            14'd10914 : begin out <= 64'b0001101111001010001010101000000010101011010001001010011101111011; end
            14'd10915 : begin out <= 64'b1010100100110110001010111110001100101000000111011010010001110101; end
            14'd10916 : begin out <= 64'b1001110000000100101010011101101100100111111001110010010100110010; end
            14'd10917 : begin out <= 64'b0010100111010001101001011111011010101001001011000010100110011000; end
            14'd10918 : begin out <= 64'b0000110111011010000110100110110000100111111000110010101011110110; end
            14'd10919 : begin out <= 64'b1010101100010000101010001101000100100111110101000010100011110001; end
            14'd10920 : begin out <= 64'b0010100011100100001010100001011010100111010001101010010000111000; end
            14'd10921 : begin out <= 64'b0001101110101001001010010100001000010110101101011010011001010000; end
            14'd10922 : begin out <= 64'b0010011001010111001010101100101000100100001110001010001100111001; end
            14'd10923 : begin out <= 64'b1010010110110111001010000101100110101011100101001010000100110000; end
            14'd10924 : begin out <= 64'b1010100110001111101010001111011010011111011111110010011001001011; end
            14'd10925 : begin out <= 64'b0010101111101001000111000010000100101011001011010010000111100011; end
            14'd10926 : begin out <= 64'b1010010111001111001000100001001110011111100100001010010001010010; end
            14'd10927 : begin out <= 64'b1010010100000000101010011011011010101000101001100010010011011000; end
            14'd10928 : begin out <= 64'b0010101100000000101010001100011100100111001101000000110000010010; end
            14'd10929 : begin out <= 64'b0010011011000100001010110001110000101001100011101010101101100010; end
            14'd10930 : begin out <= 64'b1010100110011101001010101011110110100000011100011010001110001111; end
            14'd10931 : begin out <= 64'b1010011110010101001010101110101100101011011000011010100011100001; end
            14'd10932 : begin out <= 64'b1010101110110010001010110111100100101010101011000010011100000100; end
            14'd10933 : begin out <= 64'b1010010010000111001001110111010000101000110001010001011111100010; end
            14'd10934 : begin out <= 64'b0010100010001101001001110110111010100001011110000010100110100010; end
            14'd10935 : begin out <= 64'b0001101110111000101010110111100000100100010000111001110011010000; end
            14'd10936 : begin out <= 64'b1010001110011101101001001000101000100110010101110010011010001100; end
            14'd10937 : begin out <= 64'b0010000010100111001010010011101000101000100110000010101111001000; end
            14'd10938 : begin out <= 64'b1010010010000011001010100110001010101010101110010010100101001100; end
            14'd10939 : begin out <= 64'b0001110100001000101001111011011100100010100101001001100000000000; end
            14'd10940 : begin out <= 64'b1010010011011100100111011011000100100101100011111010100001110100; end
            14'd10941 : begin out <= 64'b0010101000001101101001110100100110100101011001010010100011001110; end
            14'd10942 : begin out <= 64'b1010101101000011001010110100000100011011010110101010100000110011; end
            14'd10943 : begin out <= 64'b0010100111100011101010101100011010100110000001010010101111110111; end
            14'd10944 : begin out <= 64'b0010101011110011100110000101000000100000010110101010101110011000; end
            14'd10945 : begin out <= 64'b1010011110001111101001000111001110101001110100001010011101001111; end
            14'd10946 : begin out <= 64'b0010101010010101101001000001000110100010101011000001110011001100; end
            14'd10947 : begin out <= 64'b0001100100101110101010010101010010100110101010001010101001011110; end
            14'd10948 : begin out <= 64'b0010011000111011001001010010100100011110101000101010011011000110; end
            14'd10949 : begin out <= 64'b1010101011001000001001111101100110100010001001010010101110011110; end
            14'd10950 : begin out <= 64'b1010001111011001001010100000101100011001001110100010101111011101; end
            14'd10951 : begin out <= 64'b0010100000111011001010110100001110100001010110101010100111001000; end
            14'd10952 : begin out <= 64'b0010100000100011101001000000011010100110111110110010010110100010; end
            14'd10953 : begin out <= 64'b0001110010000111101001011001100110100100001011110010011110001010; end
            14'd10954 : begin out <= 64'b1001100111000111100111001000110100100000111001100010011011110000; end
            14'd10955 : begin out <= 64'b0010101001100100101010000010110100101001110000000010010001001110; end
            14'd10956 : begin out <= 64'b0010010111000000001001100101000100101001100001000010100001110111; end
            14'd10957 : begin out <= 64'b1001101001111011001010011111101010101001000101110010010111100000; end
            14'd10958 : begin out <= 64'b0010010010001000100110100101001010101010101010101010101010111010; end
            14'd10959 : begin out <= 64'b1010100000111001101001110010111000100100001101100010100010100001; end
            14'd10960 : begin out <= 64'b0010010111101011001010101111111110011100110010010010011111101001; end
            14'd10961 : begin out <= 64'b1010000110011011101000001111100000101011000101111001100110001011; end
            14'd10962 : begin out <= 64'b0001110000000110101000111001000110100001001000001000101101110001; end
            14'd10963 : begin out <= 64'b1010000000011110001001101111111110101011011010111010100011010101; end
            14'd10964 : begin out <= 64'b1010101000011000101001000101011110011000011100100001010000001011; end
            14'd10965 : begin out <= 64'b1010011000011010101001111111000000101000011100101010010011011101; end
            14'd10966 : begin out <= 64'b0010100000100111001010011011111100101010111001110001111100111101; end
            14'd10967 : begin out <= 64'b1010010100001100100111110110001110011110011110100010011111110100; end
            14'd10968 : begin out <= 64'b1000010001111001100111111001100010100100000110001010010100000011; end
            14'd10969 : begin out <= 64'b0001110011001001001010101011001010100100110011101010001111100011; end
            14'd10970 : begin out <= 64'b1010101100110110001010010110101110100111101111110010011010011001; end
            14'd10971 : begin out <= 64'b1010100111100010101001101111001110100110010110101010100100000100; end
            14'd10972 : begin out <= 64'b1010010111011011001010100001101100101010011111011010000011100000; end
            14'd10973 : begin out <= 64'b0010011110110001101010110000001110011110000100001010010100101011; end
            14'd10974 : begin out <= 64'b1010100000111101101010100011001010100001001010000010101100001010; end
            14'd10975 : begin out <= 64'b1010100110000011001000011100011000100001001111100010101111011111; end
            14'd10976 : begin out <= 64'b1010010011000100001010010110000000100111010110011010011001111110; end
            14'd10977 : begin out <= 64'b0010010111011011101010001000001100100010011110010010101010000001; end
            14'd10978 : begin out <= 64'b1001100101100100101010100111101010010101111001111010000001001101; end
            14'd10979 : begin out <= 64'b0010100110110101101010110111000010100111100011001010000001001100; end
            14'd10980 : begin out <= 64'b1010100001111000001010100000001100101011010101111010101011101110; end
            14'd10981 : begin out <= 64'b0010101000000011000110001011010000101010111100100010000110101110; end
            14'd10982 : begin out <= 64'b0010011100110111001010000001100000010111110100100001110100100100; end
            14'd10983 : begin out <= 64'b1010100101011001001001000101001110100111100010011010011010101001; end
            14'd10984 : begin out <= 64'b1010101001001101001010010100001010100010100111001010000011000100; end
            14'd10985 : begin out <= 64'b1010011000111110001010110110111000100111010101000001011100010010; end
            14'd10986 : begin out <= 64'b1001010011100101001010110110001000101001010101111010001000111001; end
            14'd10987 : begin out <= 64'b0001110001100100001000100010010100100010010010111010101110010010; end
            14'd10988 : begin out <= 64'b0001100110011000101010111011000010100011111100110010101000001011; end
            14'd10989 : begin out <= 64'b1010011010110101001001100010011010011010111000011010010110010101; end
            14'd10990 : begin out <= 64'b1010011010001001000100110110101100100100010101100010010010110101; end
            14'd10991 : begin out <= 64'b1000101110101001101010000101111110101011101100111001101011110011; end
            14'd10992 : begin out <= 64'b1010100000110011100111001000101000100101010110101001110111010110; end
            14'd10993 : begin out <= 64'b1010011110001001001000010101101100101011101101001010100011001111; end
            14'd10994 : begin out <= 64'b0010010100100110001010100111111000011110010111110010101001111100; end
            14'd10995 : begin out <= 64'b0010011111101000001010111110000010011110011100001010101010011101; end
            14'd10996 : begin out <= 64'b0010010101111000001010111101111000101011100001000010100101000100; end
            14'd10997 : begin out <= 64'b1010011010010100101010100010010100100100000000111010000100101001; end
            14'd10998 : begin out <= 64'b0010100010000100000101000001111100100011101001000001111110011010; end
            14'd10999 : begin out <= 64'b1010100011000101000111010000110100101011101101110010101110100100; end
            14'd11000 : begin out <= 64'b1010101110111011101001111001001110100101000001010001101111111110; end
            14'd11001 : begin out <= 64'b1001101110101111001001010001111000101000010100100010101010011010; end
            14'd11002 : begin out <= 64'b0010101010110110001001010100001110100100011010000010101000000110; end
            14'd11003 : begin out <= 64'b1010010101110101001010110100010110101010000101001001100101001110; end
            14'd11004 : begin out <= 64'b1010011001111111101010110101111110100010110100111010101101110111; end
            14'd11005 : begin out <= 64'b1001001001111100100101010101000110100001100011010010100100000011; end
            14'd11006 : begin out <= 64'b1010000111010011001010100110101110100001111011000010000111111011; end
            14'd11007 : begin out <= 64'b0010010011001110101010000110001100100101111001110010101001001110; end
            14'd11008 : begin out <= 64'b0010010011010001101010000100001110101010111111111001101110110001; end
            14'd11009 : begin out <= 64'b1010100111110101001001011011111010100111001101001010011010100101; end
            14'd11010 : begin out <= 64'b0010011111110011001001000010010110011111100101101010011011101100; end
            14'd11011 : begin out <= 64'b0001011001000001001000000011001110011010101010100010001110000000; end
            14'd11012 : begin out <= 64'b0010011111001011101010011100001100101011111001010010101101000011; end
            14'd11013 : begin out <= 64'b1010101001101111001010000001010000101000100000010010010010000111; end
            14'd11014 : begin out <= 64'b1010101011011011001010101010111100101010100100111010101000101001; end
            14'd11015 : begin out <= 64'b0010001100000111001010100001010100100001100100000010101000110101; end
            14'd11016 : begin out <= 64'b1010101110011100001000111111000110100110111101011010001010000001; end
            14'd11017 : begin out <= 64'b1010011101001011001010100111110110100000100100100010011010011110; end
            14'd11018 : begin out <= 64'b1010100101100100001010011000111000100111011110001010101011111010; end
            14'd11019 : begin out <= 64'b0010101101011001001010010000110000100101001110001010100111011000; end
            14'd11020 : begin out <= 64'b1010011011010000101001100110111110101010110011000010100011100011; end
            14'd11021 : begin out <= 64'b0010100100010000001001000101001000101000000100111010100010111100; end
            14'd11022 : begin out <= 64'b0000000001100000101010111111001100101010110011100010010110001111; end
            14'd11023 : begin out <= 64'b0010011001110111001010010011010000101011100101000010100000010110; end
            14'd11024 : begin out <= 64'b1010100101100000001010000101011100101010000100100010100010111001; end
            14'd11025 : begin out <= 64'b1010011000011001101001111101110010101000110100011010101110001100; end
            14'd11026 : begin out <= 64'b0010010110110001001010011110100100100010001101111010000111101010; end
            14'd11027 : begin out <= 64'b0010101100100001101010000010111010011110110000100010100010100100; end
            14'd11028 : begin out <= 64'b0010100110110010101001111111011100101000001001100001111111101110; end
            14'd11029 : begin out <= 64'b1001000010010011001001110100011100101001011011011010000100111001; end
            14'd11030 : begin out <= 64'b0010011101011010100110101011011010100111001110000010100101101011; end
            14'd11031 : begin out <= 64'b0001010000111010101001110101101000101001110010001010010111111010; end
            14'd11032 : begin out <= 64'b1010010101011111101010100101111010101001001010001001111100010000; end
            14'd11033 : begin out <= 64'b0010011000000111101000100101101110100001000110110010011101010011; end
            14'd11034 : begin out <= 64'b0010100100100101101000001001000000100110010101001010100011011110; end
            14'd11035 : begin out <= 64'b1001100111110111101001010001011000100110100001000010101111011011; end
            14'd11036 : begin out <= 64'b1010011111111011000111001010001110101001001000000010100010011000; end
            14'd11037 : begin out <= 64'b1010101000010001001000010100110110101000101101110010100110101100; end
            14'd11038 : begin out <= 64'b1010100110001101101010011100101100101011111011001010100111011111; end
            14'd11039 : begin out <= 64'b1010101111001110001010111000000100101010000001111010010001011001; end
            14'd11040 : begin out <= 64'b0010011001011010101010001100001000101010001000110010001010110001; end
            14'd11041 : begin out <= 64'b1010001100011011100101010110000000101011000100100010010000111101; end
            14'd11042 : begin out <= 64'b1010100001000101001001111111111100100001001000010010101000110011; end
            14'd11043 : begin out <= 64'b1010010111101011001010000011010010101000001101101010011011111111; end
            14'd11044 : begin out <= 64'b1010100110110000001001100011111010100111100101011010001001111110; end
            14'd11045 : begin out <= 64'b1010000010010011001010100100111010101001101000101010101110010000; end
            14'd11046 : begin out <= 64'b1010101000100010001000100110111000011101011100000010100001100011; end
            14'd11047 : begin out <= 64'b1010100001010011001001011101000010101001000011011010101000100000; end
            14'd11048 : begin out <= 64'b1010100100011001101001000011101100100100100111101010100111110110; end
            14'd11049 : begin out <= 64'b1010001110101111101001001010100100100001000101001010011101010100; end
            14'd11050 : begin out <= 64'b0010101000010011100110100011011000101001100100110001000111100110; end
            14'd11051 : begin out <= 64'b0001010001011111101010101000011110100001011101000010100001101100; end
            14'd11052 : begin out <= 64'b1010100010010000101000101101110000101011011100111010010010000010; end
            14'd11053 : begin out <= 64'b1010101001011101000000000111111000100111110000111010000011111010; end
            14'd11054 : begin out <= 64'b0010010010001000101010010000100000101010111011111001110000000100; end
            14'd11055 : begin out <= 64'b1010101011001010001010111011110100101010010010101010101101100010; end
            14'd11056 : begin out <= 64'b0010100000010001000111010001010110011110100101000010101010010101; end
            14'd11057 : begin out <= 64'b0010100111001110001000110101100100011110001101101010100111000011; end
            14'd11058 : begin out <= 64'b0010101001110110101010100000111100101000000101100010101000110010; end
            14'd11059 : begin out <= 64'b0010011000111000101010001111010100101010110001000010010010001100; end
            14'd11060 : begin out <= 64'b0010001101111110101010101100010010101001000110000001111101001101; end
            14'd11061 : begin out <= 64'b0010101100101011101001111111110010011111000110110010101001000000; end
            14'd11062 : begin out <= 64'b0001101000101111100111100010101000100111001010010010011010100111; end
            14'd11063 : begin out <= 64'b0010110000000001001010110110110100100010110010100010100000111111; end
            14'd11064 : begin out <= 64'b0010011100000001100111010000100110101001011111101001111111111010; end
            14'd11065 : begin out <= 64'b1010011101000101001010100011100000101000100110100010101100111100; end
            14'd11066 : begin out <= 64'b0010010110000011101001111101010010101000111110110010100110000111; end
            14'd11067 : begin out <= 64'b0001111111101101001010111110000000101010001001101010010100010010; end
            14'd11068 : begin out <= 64'b1001100011101100001010110100110110101001101010101001100100011101; end
            14'd11069 : begin out <= 64'b0010100111011010101001000111111100101001000101101010010000011011; end
            14'd11070 : begin out <= 64'b0010100011010100001010100111000100100111001101000010010010010011; end
            14'd11071 : begin out <= 64'b1001111110101111001001001000010110001101000000001010010111111010; end
            14'd11072 : begin out <= 64'b1010101011110010001001110010101110101010000110011001110100110100; end
            14'd11073 : begin out <= 64'b1001010011101101001001000111000010101011010000101001001110001111; end
            14'd11074 : begin out <= 64'b0010011001000100101001110100000110101000110110010010000001011111; end
            14'd11075 : begin out <= 64'b1001100011001001101010001110010010100011110111110010100110101100; end
            14'd11076 : begin out <= 64'b1010001110100000101001100110000010101010001101111010101100011111; end
            14'd11077 : begin out <= 64'b0010101001101101000110101111011100100000010110111010010111011001; end
            14'd11078 : begin out <= 64'b0010010010010001001010000110111110101011010001001010001100100110; end
            14'd11079 : begin out <= 64'b0010010000010000101001111010101000101000000011011001110000100010; end
            14'd11080 : begin out <= 64'b1010000011101001100111001000001000101000111100111010000011110110; end
            14'd11081 : begin out <= 64'b0010110000010010001010001000111010100111101101000010101101110101; end
            14'd11082 : begin out <= 64'b0001111011010010101001101011110110011100000001111010000101000110; end
            14'd11083 : begin out <= 64'b1010011110011110101010010011001110011110001001000010100100011101; end
            14'd11084 : begin out <= 64'b0010010010010010101010000011111110011011100101011010000001111100; end
            14'd11085 : begin out <= 64'b0010100110100010001010001001001110101001011100001010101110001110; end
            14'd11086 : begin out <= 64'b0010011100101111001010001101001000101001010010100010011101101110; end
            14'd11087 : begin out <= 64'b0010100010100000001001010001110010101001001101011010010100011011; end
            14'd11088 : begin out <= 64'b0010101110011010000111001111010000101011101110100010000101100000; end
            14'd11089 : begin out <= 64'b0010011001100000001001101101100100101000111001110010101000101011; end
            14'd11090 : begin out <= 64'b1010100011101111001010011010010110101001111100010010010000011010; end
            14'd11091 : begin out <= 64'b1010100010100111001001111000100100101010110111011010000000000010; end
            14'd11092 : begin out <= 64'b1010011110101001100110010001100100100000110111110010101010101010; end
            14'd11093 : begin out <= 64'b1010101011100110001001011101000000011110110111110010010010101001; end
            14'd11094 : begin out <= 64'b0001110100000010101010010010011110101011101000011010101111100000; end
            14'd11095 : begin out <= 64'b1010000101011111101001011101011010101000111011101010101000111011; end
            14'd11096 : begin out <= 64'b1010100101001001001010001001100110101000101101011010010010000111; end
            14'd11097 : begin out <= 64'b0010000010101111001010000000100110101000100000010010011000001000; end
            14'd11098 : begin out <= 64'b1010100101011010001010001111110110100100011101111001110010111100; end
            14'd11099 : begin out <= 64'b1010000001010101001010011010001010101011100100010010000111011001; end
            14'd11100 : begin out <= 64'b1010011001000110101000001101101100011011101010010010100111110000; end
            14'd11101 : begin out <= 64'b0010011011110000101000110000011000101010001111011010011010111110; end
            14'd11102 : begin out <= 64'b0010000010111111101000110011001010101010111011010010100100110101; end
            14'd11103 : begin out <= 64'b0010010000101111001010110101101000100000101010001010101101101110; end
            14'd11104 : begin out <= 64'b0010011111101001001010100000001010101011011111101001100110000000; end
            14'd11105 : begin out <= 64'b0010101100111010101010010100101010100111100111111010011100000011; end
            14'd11106 : begin out <= 64'b1010100001110100101001011111000100101010010110001010101010110111; end
            14'd11107 : begin out <= 64'b1001100111001011101010010100000010100111111100101010101101101000; end
            14'd11108 : begin out <= 64'b1010010111011011001010100100001000101000010110011010100101010110; end
            14'd11109 : begin out <= 64'b0001010101110011101001011000010010101010001010100001111000011010; end
            14'd11110 : begin out <= 64'b0001110010011011101010000110100000100001100001101010101000000110; end
            14'd11111 : begin out <= 64'b0001011010000000101010010001101010101011010110001010100111100101; end
            14'd11112 : begin out <= 64'b0010000000000100101001001100011010001100000101100010100011010010; end
            14'd11113 : begin out <= 64'b0010011100111110101010100101010110011000000000110010101100000101; end
            14'd11114 : begin out <= 64'b0010100010100000001001010011010110101011110100100001111110000011; end
            14'd11115 : begin out <= 64'b1010011110110000101010111000100110101010001111101010100101010110; end
            14'd11116 : begin out <= 64'b1010101001010100101010001110010110101011100001000010100000111001; end
            14'd11117 : begin out <= 64'b0010100001110001101010100001100110101000000101011010100111101010; end
            14'd11118 : begin out <= 64'b1010010000001010001000000000110010100101000010011010011101101100; end
            14'd11119 : begin out <= 64'b1010010011000011001010000111010100101011011111100010101011001001; end
            14'd11120 : begin out <= 64'b1001011101100011001010010001101000011111010111100010000110011111; end
            14'd11121 : begin out <= 64'b0001100111101111001010101010111100101011101000101010100100000000; end
            14'd11122 : begin out <= 64'b1001110101001110100110011011011110100101111110111010010001110100; end
            14'd11123 : begin out <= 64'b1010100001100101101001110010010000100011100100010010011010111010; end
            14'd11124 : begin out <= 64'b0010101110000111001001110111001100011100010011000010000011001001; end
            14'd11125 : begin out <= 64'b0010100111000111001010000101010000101001110011000010101010111101; end
            14'd11126 : begin out <= 64'b1010101000101001101010010001001010010000000101110010101001010101; end
            14'd11127 : begin out <= 64'b1010000100100011001000011001110000100110011001011010001110101101; end
            14'd11128 : begin out <= 64'b0001001000100010000101000100000010101001010111001010011011001011; end
            14'd11129 : begin out <= 64'b1010011111100000101001111111000100101001000000000010010101011100; end
            14'd11130 : begin out <= 64'b1010100100100000001000110101000000100000001100110010100111000010; end
            14'd11131 : begin out <= 64'b1010101111110010101010011000101100101011010011011010001011111110; end
            14'd11132 : begin out <= 64'b0010101001000001101010010001101010100100010101000010101001000110; end
            14'd11133 : begin out <= 64'b0001110000111001001001010000001000100110000001001010010100110110; end
            14'd11134 : begin out <= 64'b0010100011001010101001011101000110101001010001001010101110101010; end
            14'd11135 : begin out <= 64'b0001011101100101100111010101000100101000101111001010011011010010; end
            14'd11136 : begin out <= 64'b1010101000111011001001001000001110101001001011111001101111111110; end
            14'd11137 : begin out <= 64'b0010101011010110001010101111111000100101101000010010011010111101; end
            14'd11138 : begin out <= 64'b0010101010010000000110010011101010100101111011010010101100000100; end
            14'd11139 : begin out <= 64'b0010101110011011101010011011101000100100111000110010010010111010; end
            14'd11140 : begin out <= 64'b1010000101010001001010111000010100101011110001001010101110111011; end
            14'd11141 : begin out <= 64'b1010100011100101101000110001101000100110001010100010000001001001; end
            14'd11142 : begin out <= 64'b0010100100111011000111011101010010101010111100110010010001110010; end
            14'd11143 : begin out <= 64'b0010011001001000101000111011001110100110000010000010101110101110; end
            14'd11144 : begin out <= 64'b0010101111010010001001011101100000101001111000100010010000011101; end
            14'd11145 : begin out <= 64'b0010011110111110001001000010111100101001010110010010101000111011; end
            14'd11146 : begin out <= 64'b0010101001100011001001101100010010101011111110110010100001100001; end
            14'd11147 : begin out <= 64'b1010101101100100001001011011010110101011000100000010100000011110; end
            14'd11148 : begin out <= 64'b0010100011011110101001000111001110101000110110000010101011110001; end
            14'd11149 : begin out <= 64'b0010100101101111001001111100101100101010111101110010101011001100; end
            14'd11150 : begin out <= 64'b0010011010000111001000110110000000100000011100110010101011001011; end
            14'd11151 : begin out <= 64'b0010100011001110001001000000010000100101101010011010100101111000; end
            14'd11152 : begin out <= 64'b0010100011010111100111000001010010100110101001111010010100001101; end
            14'd11153 : begin out <= 64'b0010101100100010001010001001000010100101110000100010011100000000; end
            14'd11154 : begin out <= 64'b1010101001010101101010101011100100100000001010011010011100001001; end
            14'd11155 : begin out <= 64'b1010100100000010101001110110100010101010110010111010011100000011; end
            14'd11156 : begin out <= 64'b0001100000001101101010101010010110010100010000100010100011001101; end
            14'd11157 : begin out <= 64'b0000100000100011001001110101111010101001000101000010110000010000; end
            14'd11158 : begin out <= 64'b0010100101001111101010010101000100010111101000110010101011101010; end
            14'd11159 : begin out <= 64'b1010010010111001001001100001010010101010100110101010010111010100; end
            14'd11160 : begin out <= 64'b1010001101000111001010011001110000011111111101101010100011110000; end
            14'd11161 : begin out <= 64'b0010011111101000101001101001001110101011101010111010100011001101; end
            14'd11162 : begin out <= 64'b1001100110101001101010011010010110100000100111111010101010110000; end
            14'd11163 : begin out <= 64'b1010101100001010100111111001000000101011000011101010010000010000; end
            14'd11164 : begin out <= 64'b0010101001011010101010000001111010100000010110011010000000001101; end
            14'd11165 : begin out <= 64'b0010100110011001101010110011011110100100111001100010100111011110; end
            14'd11166 : begin out <= 64'b0010101010010010001000001000000110101000001010100010011001101100; end
            14'd11167 : begin out <= 64'b1010101010000111100101011111100100100110111001011010101011001101; end
            14'd11168 : begin out <= 64'b1001110101111010101001100110010100101000001011000010100010000100; end
            14'd11169 : begin out <= 64'b0010100001111010001010001011100000101000110000111010001100010111; end
            14'd11170 : begin out <= 64'b0010000100111100100110010001100100100111111110010010100011000101; end
            14'd11171 : begin out <= 64'b1010010001001000001010101111010100101011101010110010000111110010; end
            14'd11172 : begin out <= 64'b1010101010110101001010010101101000011011000100011010001110101000; end
            14'd11173 : begin out <= 64'b1010011000010110001010000000010000101011011100110001111011111111; end
            14'd11174 : begin out <= 64'b1010100000100001101001101010111100101000001010110010100110011011; end
            14'd11175 : begin out <= 64'b0010011110110101000110011110001000101011011010100010100010110100; end
            14'd11176 : begin out <= 64'b0010001001111010101001010010100010101010100001000010011110101010; end
            14'd11177 : begin out <= 64'b1001011100001101001010000110010010101011011000101010011110010101; end
            14'd11178 : begin out <= 64'b0010101010010010101000011111001010011010100101100010101011010111; end
            14'd11179 : begin out <= 64'b0001111011111000101010100001111110101001001101100010100010010101; end
            14'd11180 : begin out <= 64'b1001110101011110101010101011001000100101000100011010101001010000; end
            14'd11181 : begin out <= 64'b1010101010000101000100111011111000100010011111001010101001111111; end
            14'd11182 : begin out <= 64'b1001101001000100101010111001100010101001100011011010001100000011; end
            14'd11183 : begin out <= 64'b0010100101100110001010010011011000101000011110111010101101111101; end
            14'd11184 : begin out <= 64'b0010100101011100101010101101001010100000001000101010100001001000; end
            14'd11185 : begin out <= 64'b1001101001100111001010000000110100101000000000011010010111101000; end
            14'd11186 : begin out <= 64'b1010000100111011101001101001100000101000100111011010100000101101; end
            14'd11187 : begin out <= 64'b0010011001001111101010001011110110101011101001101010000000011011; end
            14'd11188 : begin out <= 64'b0010101000010111001000101101010100100110110101001010001010101100; end
            14'd11189 : begin out <= 64'b0010100101001011101010111011011100101001010000000010010010111110; end
            14'd11190 : begin out <= 64'b0001111100101011001010100110001100101000111000101010010101011111; end
            14'd11191 : begin out <= 64'b0010011001101101101010001111011010100100100001010010101011011001; end
            14'd11192 : begin out <= 64'b0001110000110100001001110110111000101011011101100010100100001111; end
            14'd11193 : begin out <= 64'b0010100111100110101001001100010100100110100111001010010011100101; end
            14'd11194 : begin out <= 64'b1010010101011011000111101010101110101011110100101010100100111100; end
            14'd11195 : begin out <= 64'b0010110000110001001001011100001110010011111111101001111011101011; end
            14'd11196 : begin out <= 64'b1010101100000001001000101110000010011110110101101010101111101111; end
            14'd11197 : begin out <= 64'b1010000110101100001010011110111110100110110000010010101100011001; end
            14'd11198 : begin out <= 64'b0010010000000110101010111101001000100010001111111010010010100010; end
            14'd11199 : begin out <= 64'b0010100111101101101000110001100010100101001111110010001111001100; end
            14'd11200 : begin out <= 64'b0010110000111100001001010001001110101001101010000010010000001101; end
            14'd11201 : begin out <= 64'b0010010011101110001001100001100010101011011000100010011110111110; end
            14'd11202 : begin out <= 64'b0010101010101010101010101001011000100000011101010010101101010010; end
            14'd11203 : begin out <= 64'b1010001010001111101001110011010100101011111001000010011100100110; end
            14'd11204 : begin out <= 64'b1010010111010110001010100101111000100100111110101010010010000100; end
            14'd11205 : begin out <= 64'b1010100001001101001010000111000010011011101000100001110100010010; end
            14'd11206 : begin out <= 64'b1010110000001110101001010011100100100110101100101010101111101100; end
            14'd11207 : begin out <= 64'b0010010010101101001010000110100000101001110011000010100101111011; end
            14'd11208 : begin out <= 64'b1010000101011010101010100101011010100101000100010010100101100100; end
            14'd11209 : begin out <= 64'b1010001000111001001001100011111000100101010001001010100101011100; end
            14'd11210 : begin out <= 64'b0010101101101111001010010011010010100101001010000010101011011100; end
            14'd11211 : begin out <= 64'b0010011101100001001010101001110010101011101110111001101101001001; end
            14'd11212 : begin out <= 64'b1010011110110001101010111001111010101010010111100010100011100101; end
            14'd11213 : begin out <= 64'b1010101110010011101010101111010000100011011101000010101010101111; end
            14'd11214 : begin out <= 64'b1010100011101011101010000110100100011101111110011010101110100111; end
            14'd11215 : begin out <= 64'b0010010000000110001010001110100110100101101011101010101011000000; end
            14'd11216 : begin out <= 64'b1010100010000000101010111101011110100110000101101010011111011110; end
            14'd11217 : begin out <= 64'b0010010101110100001010010011010110100111110001000010101110010101; end
            14'd11218 : begin out <= 64'b0010101110000001101010000110000100101010101001000010101000001110; end
            14'd11219 : begin out <= 64'b1010010010111101101010000110000000101010001010011010001000100111; end
            14'd11220 : begin out <= 64'b0010001111010110000111001111101100100100101010110010101111011011; end
            14'd11221 : begin out <= 64'b1001101010011100001001010100101110100101100000100010000110101110; end
            14'd11222 : begin out <= 64'b0010001010010111101010111010001110101010100000000010100010101001; end
            14'd11223 : begin out <= 64'b0010100010010111001010111001110100101000100100101010100010101010; end
            14'd11224 : begin out <= 64'b1010100011000000000111011000010100101011011100111010100001111010; end
            14'd11225 : begin out <= 64'b0001110100111101101010100111011100101100001110111010100100100011; end
            14'd11226 : begin out <= 64'b0010011010011101001010110100010010101010101110101010100110110100; end
            14'd11227 : begin out <= 64'b1010001111100100001010101101101100101001000010010001011010011001; end
            14'd11228 : begin out <= 64'b0001111011110110101001100101100010101001101010011010010101101101; end
            14'd11229 : begin out <= 64'b1010001000111010001010111001100100101011110001100010100101001110; end
            14'd11230 : begin out <= 64'b0010100101101011001010011010100100101000110011101010101001011011; end
            14'd11231 : begin out <= 64'b1010110001111100101010110001011110101000010011001001011110100100; end
            14'd11232 : begin out <= 64'b1010110000100000000111100110101100100100111001010010010101011010; end
            14'd11233 : begin out <= 64'b0010010010000011101010000110101100101010000101100010101101101001; end
            14'd11234 : begin out <= 64'b1001101010000110100110000111101000101001101111100010100111100100; end
            14'd11235 : begin out <= 64'b0010100001100010001001011101101110100001100110000010011000110010; end
            14'd11236 : begin out <= 64'b0010100110001011000100111000011100101010010111111010010000000101; end
            14'd11237 : begin out <= 64'b1010101000111101101001111010011000100011111111010010010101011100; end
            14'd11238 : begin out <= 64'b0010010100100011101010000101111110100101100101101010010110101011; end
            14'd11239 : begin out <= 64'b0010101000111000001010000000101100100111101100111010101111101000; end
            14'd11240 : begin out <= 64'b1010101010010000101001100001110100101010010101000010000011010110; end
            14'd11241 : begin out <= 64'b1010100111010110001010110011101010100010010011100010101110010000; end
            14'd11242 : begin out <= 64'b1010101111001000001010111100101100101000111011010010100110000100; end
            14'd11243 : begin out <= 64'b1010000110001110101000010010101000101010000010000010101001001101; end
            14'd11244 : begin out <= 64'b1010101101110110001010011001010110101000010111010010100100001011; end
            14'd11245 : begin out <= 64'b0010011000001111101000100101001000100100010011011010011110100100; end
            14'd11246 : begin out <= 64'b0010100110101111101010111001101100100101111111111010100110101100; end
            14'd11247 : begin out <= 64'b0010101011011111101010110101111100100100110000000010100100001110; end
            14'd11248 : begin out <= 64'b0010101000000110101010010000100000100110100101001010101010100011; end
            14'd11249 : begin out <= 64'b1010100111100001001000100111011000100110101010110010100100010101; end
            14'd11250 : begin out <= 64'b0010011010100011100110010110010110100111011100101010100000011010; end
            14'd11251 : begin out <= 64'b0010100100110100000110111110100100100011110111001010101111111101; end
            14'd11252 : begin out <= 64'b0010101111101001001010101011101000100010011100000010011011011011; end
            14'd11253 : begin out <= 64'b1010101000111100101010100000000110101000110111110010100011110010; end
            14'd11254 : begin out <= 64'b0010011011011001001001110010100100100111101010110010101101010111; end
            14'd11255 : begin out <= 64'b1010100010011100001010000110001010101011000101110010011001101110; end
            14'd11256 : begin out <= 64'b1010100010000001001010111101111100101011000000010010011000010000; end
            14'd11257 : begin out <= 64'b1010101100001000001001011001111000101000101100100010010111110100; end
            14'd11258 : begin out <= 64'b0001100110010111001010101101010010100100000100110010100000001001; end
            14'd11259 : begin out <= 64'b0001010010110001100111111010100110101001100110011010001010101110; end
            14'd11260 : begin out <= 64'b0010001010110101001000010000111110100000000010110010101010000001; end
            14'd11261 : begin out <= 64'b0010010010001000101010001001010000101001100111010010101101001001; end
            14'd11262 : begin out <= 64'b1010101011110000001000010010001010101011100110010010100000001101; end
            14'd11263 : begin out <= 64'b0010101001110011101000111111001100101011111001010010010011101100; end
            14'd11264 : begin out <= 64'b1010100000110010101010000111100100100111111011100010100010100010; end
            14'd11265 : begin out <= 64'b0010100110010110001000101001110110101010010001011010000110000111; end
            14'd11266 : begin out <= 64'b0010011100100010101010011011001000011110010011011010011000100001; end
            14'd11267 : begin out <= 64'b1010100110000010001010111011101110101001111101100010011001110111; end
            14'd11268 : begin out <= 64'b1010101100101011001010010110111100011011100100111010001101011001; end
            14'd11269 : begin out <= 64'b1010100101011100001010100000011110101001110110111010100001110011; end
            14'd11270 : begin out <= 64'b1010010111111100101010111111100100101010111110000010101010110001; end
            14'd11271 : begin out <= 64'b0010010000000001101001011111000110101011100111100010100011001000; end
            14'd11272 : begin out <= 64'b0010010101101011001001000000110100101000100100010010100110001110; end
            14'd11273 : begin out <= 64'b0010100111100101101001100111010010100001000110011010011100011111; end
            14'd11274 : begin out <= 64'b0001100010001000101001001111100010100110111100110010101010100100; end
            14'd11275 : begin out <= 64'b1010000001000111101001100101000110100101101010001010010101000100; end
            14'd11276 : begin out <= 64'b0010010001101010101010001011101110101010110010100001001011111011; end
            14'd11277 : begin out <= 64'b1010010000011111000111110011110110101001000111111010001101010001; end
            14'd11278 : begin out <= 64'b1010100101011000001001011111011110101000110110101010011100000000; end
            14'd11279 : begin out <= 64'b0010101110100010000111100000101100101001001100100001001100001110; end
            14'd11280 : begin out <= 64'b1010011111110111101010010101011110101001101110010010101101001100; end
            14'd11281 : begin out <= 64'b1010000001000011000110111001110110101000111100110010100010010000; end
            14'd11282 : begin out <= 64'b0010010100001000101010000011100010100101010000001010100010000001; end
            14'd11283 : begin out <= 64'b1000100000100100100011100010000110101000101010101001110110000101; end
            14'd11284 : begin out <= 64'b1010101010001010001010001111000000101001011000111010101111001111; end
            14'd11285 : begin out <= 64'b1010100001100010001010111010110000101001100000010010101100100101; end
            14'd11286 : begin out <= 64'b0010010011101011101001110110001000100101001100011001110100000010; end
            14'd11287 : begin out <= 64'b1010011111111100101010101010100100101010010101000010100011110110; end
            14'd11288 : begin out <= 64'b0010011011101111001010000000001010101001001100001001011101011000; end
            14'd11289 : begin out <= 64'b0010011011001100001010011010010110100101110001011010011011001110; end
            14'd11290 : begin out <= 64'b0010011001101010001001000100111000011111001000101010101000110101; end
            14'd11291 : begin out <= 64'b0010101101111100001000111000010000100110100100101010100100000001; end
            14'd11292 : begin out <= 64'b0010100001110100101001110000011000100100010010000010100001100111; end
            14'd11293 : begin out <= 64'b0010100111011111101010010000001100100011110011111010101111000100; end
            14'd11294 : begin out <= 64'b0010100001011000001000110111001010101011011010111010101110110101; end
            14'd11295 : begin out <= 64'b0001110111011011001010011101100100011111110001111010011110110011; end
            14'd11296 : begin out <= 64'b1010011000101110101010110100101010101011010101110010011011001000; end
            14'd11297 : begin out <= 64'b0010001110100001101010000011001110100111110100001010100001000001; end
            14'd11298 : begin out <= 64'b1010100011111011100111100011101000101010110111100010011101100011; end
            14'd11299 : begin out <= 64'b0010101111011010100111000011001100100101101000011010000010101101; end
            14'd11300 : begin out <= 64'b0010010110100101001010000110110110011011010001001010011011111001; end
            14'd11301 : begin out <= 64'b0010010001111110101001111111000110100101000010101010011101110100; end
            14'd11302 : begin out <= 64'b0010011010000000101010011010011010101010010001010010101100100001; end
            14'd11303 : begin out <= 64'b0010101111110110001001011011001010100100010011101010100001100001; end
            14'd11304 : begin out <= 64'b1010100100101111101010000100010110100100110010000010100100100000; end
            14'd11305 : begin out <= 64'b0010010111000000001010010011010110100111000111110010100110110101; end
            14'd11306 : begin out <= 64'b1010100101100110101010100111110110101010111110000010100110111010; end
            14'd11307 : begin out <= 64'b0010100111100100101001000101101110100110110011110010100110011011; end
            14'd11308 : begin out <= 64'b1010100100010111001010001001010110101010110100100010010111001011; end
            14'd11309 : begin out <= 64'b1001010100011111101001110111011000100000111101000010010111001010; end
            14'd11310 : begin out <= 64'b0010011000001101001010010011110110101010110111100010101011011010; end
            14'd11311 : begin out <= 64'b0010101100100111001010010100001100100110101101000010001101000110; end
            14'd11312 : begin out <= 64'b0010101001110001000101101011101010101000100110111010011110100000; end
            14'd11313 : begin out <= 64'b0010101001100000001001100010100000100111110011011010000011011110; end
            14'd11314 : begin out <= 64'b1010101011101001101000110001000010101010011000100010011111010100; end
            14'd11315 : begin out <= 64'b1010101011111111101001111111001110100111010010100010101110011010; end
            14'd11316 : begin out <= 64'b1010001101010001101010001011101110100101001110101010101011110011; end
            14'd11317 : begin out <= 64'b1010001001000010101000111000010000101000111101110010001100010110; end
            14'd11318 : begin out <= 64'b1010100100111100101010010010100110101010000101111010010101110110; end
            14'd11319 : begin out <= 64'b1010101100111110100000001101001000100100111111100010100101100000; end
            14'd11320 : begin out <= 64'b0010101001000110001000111100110000100110110011010010100010111101; end
            14'd11321 : begin out <= 64'b1010011101001011001010001100111110100101010010011010100011111001; end
            14'd11322 : begin out <= 64'b0010100111100101101001101101011010101000101000110010000010000001; end
            14'd11323 : begin out <= 64'b1010101101011101101001000010001000100001001010001010100100110111; end
            14'd11324 : begin out <= 64'b1010101010111100000101110001001100100101101110010010101010010111; end
            14'd11325 : begin out <= 64'b1010101000001110001010101111100100100110110100001010011010010101; end
            14'd11326 : begin out <= 64'b0010011111100101101000100011100110100010001111111010101111010010; end
            14'd11327 : begin out <= 64'b0001110011010101101010011111010010100111110000110010011001100111; end
            14'd11328 : begin out <= 64'b0010000011110101101010001100011000100000011010010010100111001100; end
            14'd11329 : begin out <= 64'b0010100011011001101001101001000100100001100101010010011001000100; end
            14'd11330 : begin out <= 64'b1010011100001010000110010101001010100101100110110010101001011111; end
            14'd11331 : begin out <= 64'b0010100011010110101010001110110110101001100001111010100111010100; end
            14'd11332 : begin out <= 64'b0010100010001000101000111110011000100010101000010010100100000101; end
            14'd11333 : begin out <= 64'b0010101011101000101000111111111010010101001011110010100101111001; end
            14'd11334 : begin out <= 64'b1001100011001100101010001001110000101000010010010010011111000010; end
            14'd11335 : begin out <= 64'b0010011011010000001001110011101100100111011010010010010111100010; end
            14'd11336 : begin out <= 64'b1010100110100110101010101010000110101010110110010010101110000101; end
            14'd11337 : begin out <= 64'b0010101000001010001000101110010100101010100101011010101111011111; end
            14'd11338 : begin out <= 64'b0010100110111111100110110000011010100011110011001010011110001110; end
            14'd11339 : begin out <= 64'b1010101101110001101010101011100100100100010011011010100101111101; end
            14'd11340 : begin out <= 64'b1010000010110001001010101110100110101010010100101010100111000000; end
            14'd11341 : begin out <= 64'b0001101011110110001001110011001010100110010111010001010100111110; end
            14'd11342 : begin out <= 64'b0010100110111100101010000000000000101011110001101010101110010110; end
            14'd11343 : begin out <= 64'b0010101100011001101010111010111100011110000011011010101111010100; end
            14'd11344 : begin out <= 64'b0010101111001111001010110110111100101000001001010010010000110000; end
            14'd11345 : begin out <= 64'b1010100011010100101010100100101110101011111110011001111011000001; end
            14'd11346 : begin out <= 64'b0010000100101000100111011011001010100101111111100010101000000001; end
            14'd11347 : begin out <= 64'b0010010001111101000111111010011100101000100111011010100101101100; end
            14'd11348 : begin out <= 64'b1010100110111100101000001010110110100101100001011010000011111000; end
            14'd11349 : begin out <= 64'b1010101000100010101001110001101000101011001111001010000010111011; end
            14'd11350 : begin out <= 64'b0010101110100101101001000101100110011101111100011001111011000001; end
            14'd11351 : begin out <= 64'b0010101011010100100100000111011000101000011101101010010001011110; end
            14'd11352 : begin out <= 64'b1010101000101011101010100101010010100001000101000010100111011001; end
            14'd11353 : begin out <= 64'b0010100101110000001000000101010000101001110011000010100101011111; end
            14'd11354 : begin out <= 64'b0010101101100011100110001100110100011100000101110010010001100001; end
            14'd11355 : begin out <= 64'b1010011101101011101010111000111000100011010001001010011011000111; end
            14'd11356 : begin out <= 64'b1001010010001001101010110111011100100110100111101010100101100010; end
            14'd11357 : begin out <= 64'b0010101110101101001010000011000110101000101111001010100100100010; end
            14'd11358 : begin out <= 64'b0010100011000001001010110110100000101010001110001010011000100010; end
            14'd11359 : begin out <= 64'b1010010010111001001010101101011100011010001000100010101100001110; end
            14'd11360 : begin out <= 64'b0010010101001101001010100101001100101000110100001010100000110100; end
            14'd11361 : begin out <= 64'b1010001101011000100110110101000000100111101000101010100010001011; end
            14'd11362 : begin out <= 64'b0010011110110111001010110011101000101011110110101001111101011111; end
            14'd11363 : begin out <= 64'b0001001000000011001010100111000010100101101001110010100101110000; end
            14'd11364 : begin out <= 64'b0010101101110111101010011100011100101000011000000010101011011110; end
            14'd11365 : begin out <= 64'b1010011101111010001010110000111000011001011100001010101011111101; end
            14'd11366 : begin out <= 64'b1010101110100011000111101001100110101010101001110010011000100111; end
            14'd11367 : begin out <= 64'b0010010001000111001010100001010010100001011101000010011110111000; end
            14'd11368 : begin out <= 64'b1010100111001100101000011111001100101011011110001001100111001101; end
            14'd11369 : begin out <= 64'b0001111001100101101010110011111010101001101000010010011101110010; end
            14'd11370 : begin out <= 64'b1010100111000111101000000100101110011111110000110010100111111101; end
            14'd11371 : begin out <= 64'b1010000111110010001010000000011100010001100111101001100010100011; end
            14'd11372 : begin out <= 64'b0010011011000111001010101101001110100010110100100010001010010000; end
            14'd11373 : begin out <= 64'b0010000111010000000111001110111010100101010111110010101001010000; end
            14'd11374 : begin out <= 64'b1001100111010000001010011010100100101011101001101010101100001000; end
            14'd11375 : begin out <= 64'b0010011000001110001000010001001110100100001001010010100111101111; end
            14'd11376 : begin out <= 64'b1010011001001100001000011111111000101010110001110010100011011111; end
            14'd11377 : begin out <= 64'b0010001110010100001010011110100010100111010000110010011111110111; end
            14'd11378 : begin out <= 64'b1010010001000011101010001000101010100101110101000010101001000111; end
            14'd11379 : begin out <= 64'b1010100100000110001001111101011010100011001001110010101101010100; end
            14'd11380 : begin out <= 64'b0010100101000111101001101101100000100100101011000010011101110011; end
            14'd11381 : begin out <= 64'b0010000111010110101010000000101100100100111000000010100011111001; end
            14'd11382 : begin out <= 64'b0010001100110100101001110001011000101011000011100010101111100011; end
            14'd11383 : begin out <= 64'b0010011101011001101001000010001000100100001011111010100101101101; end
            14'd11384 : begin out <= 64'b0010101001111000101010101001001000100100101100000010011100110001; end
            14'd11385 : begin out <= 64'b0010000011111100001010001001010000100111100101101010101000110111; end
            14'd11386 : begin out <= 64'b0001110000111000101010001000011100101000100101110010100101111000; end
            14'd11387 : begin out <= 64'b0010101111010011001001110101100100100111110100010010101101011100; end
            14'd11388 : begin out <= 64'b0010010100011111001000110100010100101010110010000010100111100100; end
            14'd11389 : begin out <= 64'b1010110000010110101000011010111000101011100000101010000111111101; end
            14'd11390 : begin out <= 64'b1010101011101001101010000011110010100000111101101010100110011011; end
            14'd11391 : begin out <= 64'b1010100101100111101001010111010010001000001100100010100110010100; end
            14'd11392 : begin out <= 64'b1010011100100001101010010010010100100110100001010010101011100111; end
            14'd11393 : begin out <= 64'b0010100011001111101010011101000100100110001101001010010000111000; end
            14'd11394 : begin out <= 64'b0010001011000100101000100000100000100110110010010001111011010010; end
            14'd11395 : begin out <= 64'b0010100110000011000111100101001100100011001011111010100000101111; end
            14'd11396 : begin out <= 64'b1010101110001000101010011010001000101010000110001010101010000001; end
            14'd11397 : begin out <= 64'b1010101010100000000110000110110000100001100000011010000110000101; end
            14'd11398 : begin out <= 64'b1010100000010100001010110000010110101011111101001001110100000010; end
            14'd11399 : begin out <= 64'b1010100001111001001000110011110010101011010011111010010001101011; end
            14'd11400 : begin out <= 64'b1001001111001010001010000100001010101010110000111010100010001001; end
            14'd11401 : begin out <= 64'b0010000111101001101010001001010100101010010010100010100111000101; end
            14'd11402 : begin out <= 64'b0010010001101111101010011110011110011100010011001010100000000011; end
            14'd11403 : begin out <= 64'b1010100100000010001001011111111110101010101100100001010101110010; end
            14'd11404 : begin out <= 64'b1010100000100111101010111011100110011101110011100010010111100111; end
            14'd11405 : begin out <= 64'b0010101011110110001010110011010000100111001001101001110100100001; end
            14'd11406 : begin out <= 64'b1010100000100000101010110110001010010110010100101010100110101011; end
            14'd11407 : begin out <= 64'b0010001101110001101000011101101110100010111001001010100111000101; end
            14'd11408 : begin out <= 64'b1010100111011000001001100001011100101011011010000010100011100110; end
            14'd11409 : begin out <= 64'b1010100000100010001001001011001110011001000010011010101001101111; end
            14'd11410 : begin out <= 64'b0010101100100111001010000001011100101011001011111010101001001011; end
            14'd11411 : begin out <= 64'b1010100010110001101001011010011100101011010111000010100010010101; end
            14'd11412 : begin out <= 64'b0010100110001000001010000000110010101000010100111010000011101101; end
            14'd11413 : begin out <= 64'b1010100010000110101001110100000010011101111111100010000111011100; end
            14'd11414 : begin out <= 64'b0010101000110110101001011011000110100011010111000010100001001001; end
            14'd11415 : begin out <= 64'b1010101111110101001001101101110100101010110010010010101101001000; end
            14'd11416 : begin out <= 64'b1001011010000001000111101101100010101011110111001010100011000101; end
            14'd11417 : begin out <= 64'b0010101000110010101010111100100110100110111011001010011000010000; end
            14'd11418 : begin out <= 64'b1001101100010110000111100000001100101000110110100010001000000101; end
            14'd11419 : begin out <= 64'b0001110111010111101000110001101010100101110110111001011101100100; end
            14'd11420 : begin out <= 64'b1010100101110011101010000100100100011110010001001010011000011011; end
            14'd11421 : begin out <= 64'b1010101011000110100110100011101100101000000010101010010110101111; end
            14'd11422 : begin out <= 64'b0010100000100010001000010011001010100101110000101010101110100110; end
            14'd11423 : begin out <= 64'b0010011000110010101001010111000010101010000001010010100100001110; end
            14'd11424 : begin out <= 64'b0010100110000000100011000001110000001101111010100010100010010101; end
            14'd11425 : begin out <= 64'b1010010111101100101010110000001110100100011101111010100101101000; end
            14'd11426 : begin out <= 64'b1010100111100001101001101101110110101000000011010010011100001100; end
            14'd11427 : begin out <= 64'b0010100100011010001010101000111000101010111100011010011010011100; end
            14'd11428 : begin out <= 64'b0010100000111011101010100000011000100011000100000001111100011110; end
            14'd11429 : begin out <= 64'b0010000011001100101001010100101010100001111000110010000111010101; end
            14'd11430 : begin out <= 64'b1010001000111100001001011101001110100010110110001010010010011110; end
            14'd11431 : begin out <= 64'b0010011110010011001001001010010000101000101101100010011010010000; end
            14'd11432 : begin out <= 64'b1010010001011010001010110100110000101001111001100010101100001101; end
            14'd11433 : begin out <= 64'b1010100100000001100101110000011110100010011111110010001001011111; end
            14'd11434 : begin out <= 64'b0010000111011001100011100011010010101011101010011010000111111101; end
            14'd11435 : begin out <= 64'b0010010000110001000110001001010110011010010001011010100010110011; end
            14'd11436 : begin out <= 64'b1010000000010011001001011011100110101011111011001010101010101110; end
            14'd11437 : begin out <= 64'b0010011111011001101010110101000100100010101100111010100111001010; end
            14'd11438 : begin out <= 64'b0010001111101000101010101001000110100100110001001010011001110010; end
            14'd11439 : begin out <= 64'b1010001001110011101001110111110100100110100111111001100110111100; end
            14'd11440 : begin out <= 64'b0010101000111010101010010000101010101010101011011010100010111111; end
            14'd11441 : begin out <= 64'b0010100000011111001010010101101010101011111010001010100101001011; end
            14'd11442 : begin out <= 64'b0010011011000011100111100111100010011111111010100010011010100010; end
            14'd11443 : begin out <= 64'b0010100100010001001010011110100100101010110110011010100011111111; end
            14'd11444 : begin out <= 64'b1010010110111110101010110110000010101010000001000010011010000111; end
            14'd11445 : begin out <= 64'b0010100110011000101010001011111010101011010010100010010111001110; end
            14'd11446 : begin out <= 64'b0010101001110010001000110000111100101001011101010010010100000010; end
            14'd11447 : begin out <= 64'b1010100110111011001010101010010000100000010110100010000110110111; end
            14'd11448 : begin out <= 64'b0010110000010010001010101001001100100111110010000010000000100101; end
            14'd11449 : begin out <= 64'b0010100001101111100100100001101100101010000110011010000000001111; end
            14'd11450 : begin out <= 64'b0010100011010101101010001011000100101011110111111010100111110101; end
            14'd11451 : begin out <= 64'b1010101000100100101000001000111000101000000100110010000000010110; end
            14'd11452 : begin out <= 64'b0001101100101000100110011101111000100110011110001001110000101100; end
            14'd11453 : begin out <= 64'b1010101000110001001001000001111110101010000011101010001010010101; end
            14'd11454 : begin out <= 64'b0010011110111110001001101110110010101001100101010010010111101100; end
            14'd11455 : begin out <= 64'b1001110011011000101010111000000000101001110001011010000011011110; end
            14'd11456 : begin out <= 64'b1010101110001101101010011100100000101001101110100001101011101010; end
            14'd11457 : begin out <= 64'b0010010000101101101010101001111110101000001101101010011000010111; end
            14'd11458 : begin out <= 64'b1010011011000111101010111110000000101000110100010010011011100111; end
            14'd11459 : begin out <= 64'b1010101110001011001000100010010110101000100101101010100001001011; end
            14'd11460 : begin out <= 64'b1010100010000111101000010001010110100011101001011001101110010110; end
            14'd11461 : begin out <= 64'b0010100000100011001001000100010010100010001001101010010101111011; end
            14'd11462 : begin out <= 64'b0001011101111101001001100101001100101011110011101010011100000110; end
            14'd11463 : begin out <= 64'b0010100000011111001010111101011110100110011011000010101001110111; end
            14'd11464 : begin out <= 64'b1001001001001010101010001000010010101000110111101001110111011000; end
            14'd11465 : begin out <= 64'b1010001100101001001010101010101000101010100101001010100100110000; end
            14'd11466 : begin out <= 64'b0010100010101011101010100001001000101001010011010010010110110111; end
            14'd11467 : begin out <= 64'b0010100100000001001010110001000110011100110000110001111010001001; end
            14'd11468 : begin out <= 64'b1010001000101110001000000000000110101000100011000010101111010011; end
            14'd11469 : begin out <= 64'b1010101001001110001010000100000010101010010000101010100010100001; end
            14'd11470 : begin out <= 64'b0010100100011110101010101101101010011111100101100010000001011010; end
            14'd11471 : begin out <= 64'b1010101011010110001001011010111000100110110100000010011100010111; end
            14'd11472 : begin out <= 64'b0010100111010010000110111010101010101010110110011010101011100000; end
            14'd11473 : begin out <= 64'b1010100000100000001000011110111100101000101000011001000101000001; end
            14'd11474 : begin out <= 64'b0010011101000111101010101110001100101000100100110010101110101000; end
            14'd11475 : begin out <= 64'b0010101101101010101010000000101010100100010110111001010110111011; end
            14'd11476 : begin out <= 64'b1010100111100011101001000101100000101011010000010010100101010101; end
            14'd11477 : begin out <= 64'b0010001011010011101001000011101010100101010001101010100110001000; end
            14'd11478 : begin out <= 64'b1010101111101101000111101110010000100111111000101010100010110111; end
            14'd11479 : begin out <= 64'b1000100101101110001001100111011110101010001110000010101011001011; end
            14'd11480 : begin out <= 64'b1010101111111001100011000101000000101010111011100010101101110100; end
            14'd11481 : begin out <= 64'b1010100011110110101010011010111010100101111100100001110101001110; end
            14'd11482 : begin out <= 64'b1010000111001000101001011111101010100100001001101010101111011001; end
            14'd11483 : begin out <= 64'b1010101011101101000111101111000100100010001000100001111011001011; end
            14'd11484 : begin out <= 64'b0010101101001111101010110011010000101000111011010001100001101001; end
            14'd11485 : begin out <= 64'b1010101000011001101010011001001100100011111101100010100001111101; end
            14'd11486 : begin out <= 64'b1010101101100001101010000001110000100110110110010010101011111111; end
            14'd11487 : begin out <= 64'b1010101001100000100111000001100100101000101100101010001110101100; end
            14'd11488 : begin out <= 64'b0001101010000111101010101100100000100100010001111001001101101110; end
            14'd11489 : begin out <= 64'b1010101110001100101010011100100100100101001111010010101100010011; end
            14'd11490 : begin out <= 64'b1010101111001011100101000111010110101010010100010010100011111010; end
            14'd11491 : begin out <= 64'b1010000001101101101010101010000110100010101101101010010001101100; end
            14'd11492 : begin out <= 64'b1010101110111011100001101010001110101011010110010010100010000011; end
            14'd11493 : begin out <= 64'b1010100101000101000111100101111000101011100001100010000100000010; end
            14'd11494 : begin out <= 64'b1010101001011101101010101101001010101011111010110010100001110001; end
            14'd11495 : begin out <= 64'b1010010100100110001010111101011110101001011001101010100000111011; end
            14'd11496 : begin out <= 64'b1010101000110000100111001010101000101000110110111010011010010111; end
            14'd11497 : begin out <= 64'b0010100001000110001010111100111100001111101111010010100001010001; end
            14'd11498 : begin out <= 64'b1010001110101011001010011011101010101000011011101010010000000011; end
            14'd11499 : begin out <= 64'b1010100101010011001010111100111000101011001011000001111101000001; end
            14'd11500 : begin out <= 64'b1001111001111110101010111001001000101001011100100010010010110001; end
            14'd11501 : begin out <= 64'b1010000001000000001010010001111100101010100100101010011101110011; end
            14'd11502 : begin out <= 64'b0010100111101101001001110010010110101011100100101010100000100110; end
            14'd11503 : begin out <= 64'b1010010101100001101010001111100100101000100100101010010011101011; end
            14'd11504 : begin out <= 64'b0010000011000011001000000001001010100101100001011001110001100011; end
            14'd11505 : begin out <= 64'b1010101011101000101010000010100010100101011000010010101111010110; end
            14'd11506 : begin out <= 64'b0010101000110100001010010000011000100000110110100010101101111000; end
            14'd11507 : begin out <= 64'b0010001000110011001001011001111110100100001110000010100101110011; end
            14'd11508 : begin out <= 64'b1010010111001000001010111110101000100111110111011001100110011111; end
            14'd11509 : begin out <= 64'b0010100100100111001001110010001100100101110010101010011000011101; end
            14'd11510 : begin out <= 64'b0010101101100110001001011111001110100111010000110010010010000001; end
            14'd11511 : begin out <= 64'b0010101010011100000111010101011000101011010100000010011111011111; end
            14'd11512 : begin out <= 64'b1010011001100110001000011110100000100101110110001010000101010010; end
            14'd11513 : begin out <= 64'b1010010000010011101010101010000100101000110000001010010011001110; end
            14'd11514 : begin out <= 64'b0010101000000101101010110100011110100101110000111010101100000010; end
            14'd11515 : begin out <= 64'b1010101011101000101010111001101100101010100111111010101101010001; end
            14'd11516 : begin out <= 64'b0010101011111000001010100000000010100100000010001010100111100101; end
            14'd11517 : begin out <= 64'b1010100111000110001000000110110010100101101111101010100110100101; end
            14'd11518 : begin out <= 64'b0010101101101111001010011001101100101001110110010010100101111101; end
            14'd11519 : begin out <= 64'b0010100111111001001001011111101100101010001110010010100100110111; end
            14'd11520 : begin out <= 64'b1010011010000101000111110110001000100100001100000010100010110010; end
            14'd11521 : begin out <= 64'b0010100010100000001001010100111100011111100000111010000111110100; end
            14'd11522 : begin out <= 64'b0010100110000111101010001001010000100011110100111010010110110111; end
            14'd11523 : begin out <= 64'b1010100110100100001010111111111010010100111010111010001011110010; end
            14'd11524 : begin out <= 64'b1010100100111101101010101100011110100110100010101001101011010100; end
            14'd11525 : begin out <= 64'b0010010010010110101010010100101110100100111011101010101111010001; end
            14'd11526 : begin out <= 64'b1001111011000110101000101010000010101011100101110001110111111001; end
            14'd11527 : begin out <= 64'b1010100010000011101010111011011100011100110100111010100000001000; end
            14'd11528 : begin out <= 64'b1010100001000000101001100000111110101011101101110001110011110111; end
            14'd11529 : begin out <= 64'b1010011001101111001000111111011010100100000011111010011000001111; end
            14'd11530 : begin out <= 64'b1010011011111001000110011010100110011010111111000010100001011001; end
            14'd11531 : begin out <= 64'b0010001100100000001010000000110110100110101100101010010011110011; end
            14'd11532 : begin out <= 64'b1010011001010100101010111011010110101010110001010010011010110010; end
            14'd11533 : begin out <= 64'b1001110011101000001001000100010000101000001010010010101000111111; end
            14'd11534 : begin out <= 64'b1010101010000010001010100101001000101010101010110010100110101010; end
            14'd11535 : begin out <= 64'b0010100101101010101010001110111010100111001111101010001101110101; end
            14'd11536 : begin out <= 64'b1010011101001010001010001111110100101000001110001010010100000101; end
            14'd11537 : begin out <= 64'b0010101101001000101010110111110100101001001100010000110110000001; end
            14'd11538 : begin out <= 64'b1010010010010011101010011000011010100100111111111010000111011111; end
            14'd11539 : begin out <= 64'b0010100000010010101010000110011000100101110010001001110110011001; end
            14'd11540 : begin out <= 64'b1010100110110000101000111110011000101011111100010010101001011000; end
            14'd11541 : begin out <= 64'b0010100100000101101010111010000110101011000000101010100100011101; end
            14'd11542 : begin out <= 64'b1010011010011100101001011101110000100101100011011010001011011101; end
            14'd11543 : begin out <= 64'b0010011001111001001001101101110010011110000000111010100010010110; end
            14'd11544 : begin out <= 64'b1010010000000010101001000001011100010100011100101010101001000100; end
            14'd11545 : begin out <= 64'b0010101010110010100101010110101100100111011011110010101010001010; end
            14'd11546 : begin out <= 64'b1010100001111111001000111011010110101010010010100010000011001011; end
            14'd11547 : begin out <= 64'b0010000000000100001010011100111100100011101101100010000011010100; end
            14'd11548 : begin out <= 64'b1010000000000110001010101011111110101000110111111010011010000011; end
            14'd11549 : begin out <= 64'b0010001100001011001000010100001110101000101100100010101001110001; end
            14'd11550 : begin out <= 64'b1010011101101000101010100110010100101010010100111001011000110101; end
            14'd11551 : begin out <= 64'b1010101000010101101010001000001010101011011000010010000011111110; end
            14'd11552 : begin out <= 64'b0010100110010001101010101101001100100000000011001010100001010000; end
            14'd11553 : begin out <= 64'b1010011011101010000111110110100010101001101111010010010000111001; end
            14'd11554 : begin out <= 64'b1010011011110011001010100101110010100111010100000010101110100110; end
            14'd11555 : begin out <= 64'b0010100100000010100101001101101110101001011000110010101010101101; end
            14'd11556 : begin out <= 64'b0001111001000100101010111011011110010011101110111010001110000101; end
            14'd11557 : begin out <= 64'b0010101100101000101000000001011110100100100101111010011011101010; end
            14'd11558 : begin out <= 64'b0010100001100101001010101010000010101011001001010010000011111000; end
            14'd11559 : begin out <= 64'b1010011011011100001001001010011110101011110110011010001110000110; end
            14'd11560 : begin out <= 64'b1010011011001110001010001100001100100000100101111010011011000000; end
            14'd11561 : begin out <= 64'b1010100011110010101010101011000110011100010110110010100011000011; end
            14'd11562 : begin out <= 64'b1010000001110010101001011000011110101011110000010010101000101100; end
            14'd11563 : begin out <= 64'b0010101010101101000101001111111100101001111011110010100111100011; end
            14'd11564 : begin out <= 64'b0010101001001101000111100001011010011110011001010010100000111101; end
            14'd11565 : begin out <= 64'b1010100100110111001010010000110010011101110000000001111010110011; end
            14'd11566 : begin out <= 64'b0010101100101010001000000001101000101000010000011010000110101001; end
            14'd11567 : begin out <= 64'b1010101010010110101001110000111100101001011010110010101010011011; end
            14'd11568 : begin out <= 64'b0010101011011010001001110110111100101010011100011010101010001001; end
            14'd11569 : begin out <= 64'b0010011010000111101010010110011100101001110110110010000001111001; end
            14'd11570 : begin out <= 64'b0010010110000100101001110000111100101000101111011010010000101100; end
            14'd11571 : begin out <= 64'b1010001000111111001010001011111110100101100111001010010010100000; end
            14'd11572 : begin out <= 64'b1010100000111111101010111001101110101000011100011010000110000011; end
            14'd11573 : begin out <= 64'b1010100000000010001010111010111110101010100110000010011100001000; end
            14'd11574 : begin out <= 64'b0010010011101011101000010000100110011111010100001001111001110110; end
            14'd11575 : begin out <= 64'b0010100101111100101010000000101000011000000110100010011001010001; end
            14'd11576 : begin out <= 64'b1010011100000111000111001011000010101011011001100010100100000011; end
            14'd11577 : begin out <= 64'b0010001001110000101010111111110000101001001100111010100000101101; end
            14'd11578 : begin out <= 64'b1010010000011011001010011000111110101000111111000010011010100101; end
            14'd11579 : begin out <= 64'b0010010000001000001010110011001110101001100011001001111100101110; end
            14'd11580 : begin out <= 64'b0010101100110000101011000000000000100001110010111010101100001010; end
            14'd11581 : begin out <= 64'b1010000100111010001001010110111110101001100000001010000100110111; end
            14'd11582 : begin out <= 64'b0010100010000110001010010001111010101011101001001010011001110110; end
            14'd11583 : begin out <= 64'b0010100101011111001001101101001100011001010010100010101000000010; end
            14'd11584 : begin out <= 64'b0001111001011100001010100011111000100011100110101010010111001010; end
            14'd11585 : begin out <= 64'b1001101110001100101010011000100100101011101000011010101101000111; end
            14'd11586 : begin out <= 64'b1001100101111101101010001100010100100101000100110010100001101001; end
            14'd11587 : begin out <= 64'b1001111011101111100111011110101100101000101111111010100110000110; end
            14'd11588 : begin out <= 64'b1010100001000100001010010110110110100010100111010010011000110001; end
            14'd11589 : begin out <= 64'b0010011110010001001010100001001100100110000011101001110111011110; end
            14'd11590 : begin out <= 64'b0010011001000101101010110011101110101000110010110001100010110111; end
            14'd11591 : begin out <= 64'b0010101111100110001010111010100010101010001000101010101101010110; end
            14'd11592 : begin out <= 64'b0001011000111011001001001100100110100010100000001001011110010101; end
            14'd11593 : begin out <= 64'b0010011000011011000111000101101110011111011001111010100110100001; end
            14'd11594 : begin out <= 64'b1010011000111010101010011111011110101001010001100001101000010001; end
            14'd11595 : begin out <= 64'b0010100000011010100110010100101000101000010000010010100101100110; end
            14'd11596 : begin out <= 64'b1010000101101101100111001010111100101000011100011010010001110110; end
            14'd11597 : begin out <= 64'b0001110010111111001010100101001010011110101000101010100100110001; end
            14'd11598 : begin out <= 64'b1010011101110101101010101100100110000111111010110010010011100100; end
            14'd11599 : begin out <= 64'b0010011001010110001010011001100010101000000011111010100011100000; end
            14'd11600 : begin out <= 64'b1010010110000101001010011000011010100011100100011010011001111101; end
            14'd11601 : begin out <= 64'b1010101010001110101010111100110000101001001101011010101010000010; end
            14'd11602 : begin out <= 64'b1010101001111110100110001011111010100111100011010010101001000001; end
            14'd11603 : begin out <= 64'b1001101110001100001010001010001110011100001110111010101000011100; end
            14'd11604 : begin out <= 64'b1010000101001000001010110101100010010100101111111010011100000000; end
            14'd11605 : begin out <= 64'b0001100110010100001010011101001110100001010100110010100010010111; end
            14'd11606 : begin out <= 64'b1010011110001010100010001001111110101010111001001001110011011101; end
            14'd11607 : begin out <= 64'b0010011100011000001010110110010100101001011001100010101000010101; end
            14'd11608 : begin out <= 64'b1010101101011110001010111100110100011001101101011010101100111110; end
            14'd11609 : begin out <= 64'b0010100000001011101010010100010000100000110011010010101011110011; end
            14'd11610 : begin out <= 64'b1010010110110010001010011000011000101001001011011001111010111111; end
            14'd11611 : begin out <= 64'b1010100011101110101010111101100110101010101101000010101100110000; end
            14'd11612 : begin out <= 64'b0010101001100001101000100111111110100110100000010010110000110110; end
            14'd11613 : begin out <= 64'b1001110001001000101001000010000010100001110101011010100011110100; end
            14'd11614 : begin out <= 64'b0010101011000110001010001100110000011101110001001010100001000100; end
            14'd11615 : begin out <= 64'b0010101101110100001010000011101010100100101100100010101100101110; end
            14'd11616 : begin out <= 64'b0010010011001110001010010000000010101001010111001010100111101000; end
            14'd11617 : begin out <= 64'b0010011111001010101010011110011010101010011100100010100110010111; end
            14'd11618 : begin out <= 64'b0010101111101101001010010110101110101000011000010010101100110001; end
            14'd11619 : begin out <= 64'b1010010100101001101010101000110110101000011110100010011100010101; end
            14'd11620 : begin out <= 64'b1010100000000010101001111101000000101011011110011010101111000011; end
            14'd11621 : begin out <= 64'b1010010110011100101000000100100110101001000010001010010110010001; end
            14'd11622 : begin out <= 64'b1010101000000000000110101000001100101011011100111010101101000001; end
            14'd11623 : begin out <= 64'b0010101010101000001000100110000100100011101010100010000111011010; end
            14'd11624 : begin out <= 64'b1010101011000001001010001111000000011100001010110010000001101000; end
            14'd11625 : begin out <= 64'b1010010101010011100011111011011010100101001111110010101110010111; end
            14'd11626 : begin out <= 64'b1010010110110000101010010101101000100111001110011010000000100000; end
            14'd11627 : begin out <= 64'b0010010000010101101001000000010000100010011001111010011101101001; end
            14'd11628 : begin out <= 64'b0010101011110111001001110011011100101011100001001010011001010000; end
            14'd11629 : begin out <= 64'b0010100101010011101010111110101110100110010110100010101001111010; end
            14'd11630 : begin out <= 64'b1010011010111110001010001000000000010111010001101010011100011110; end
            14'd11631 : begin out <= 64'b1010101100101101101010001111110110101010100101101010101011010000; end
            14'd11632 : begin out <= 64'b0010011000110110001000011000001100101000000010101010100010100011; end
            14'd11633 : begin out <= 64'b1010010011101111001010111110111110101010110011100010100101101001; end
            14'd11634 : begin out <= 64'b1010010110111000101010000101000110010110011100001010101010000101; end
            14'd11635 : begin out <= 64'b1010100010000011001001100101101000101000110000111010100010001100; end
            14'd11636 : begin out <= 64'b1001001100011111100101110111001010101011110100011010100000010100; end
            14'd11637 : begin out <= 64'b1010011011011101101010101111010110100000111010100010100110100110; end
            14'd11638 : begin out <= 64'b1010101011000101001010111000010000011011111111010010011011111101; end
            14'd11639 : begin out <= 64'b0010100000001011101001110111101100101010011011110010101101010000; end
            14'd11640 : begin out <= 64'b0010001111110111101010101100111110010100110110111010100011001110; end
            14'd11641 : begin out <= 64'b0010100001100101001010001110110010100101011100111010100111001110; end
            14'd11642 : begin out <= 64'b1010010000101010101000010000010110101011110011000010110000000110; end
            14'd11643 : begin out <= 64'b1010100000101001001001000110011100100111010101100010011011101101; end
            14'd11644 : begin out <= 64'b0010100000000101101010111011111110011110001100101010101100110001; end
            14'd11645 : begin out <= 64'b0010100110111010101000101010101000101010111000100010100111011101; end
            14'd11646 : begin out <= 64'b0010001011110100000111101110110100101011010100111010101110111101; end
            14'd11647 : begin out <= 64'b0010010010111110001001100001110110011000001111111010101101110001; end
            14'd11648 : begin out <= 64'b0010010001101100001001111101100000101000010000000010000101110111; end
            14'd11649 : begin out <= 64'b1010100111110101000111110101101100101000010010110010100101011100; end
            14'd11650 : begin out <= 64'b1001100000101101101001111101110010100110111101010010011100110011; end
            14'd11651 : begin out <= 64'b0010101011110011001001111110001010100011010011011010100011100000; end
            14'd11652 : begin out <= 64'b1010101001110110100111010111000110100100010101110010101000011110; end
            14'd11653 : begin out <= 64'b1010101011101111001001011011011100101000100011101010100110110011; end
            14'd11654 : begin out <= 64'b0010001011010110101010100101110000101100001011001010100000101001; end
            14'd11655 : begin out <= 64'b1010101001101110101010100000001000101011011011011010011000110101; end
            14'd11656 : begin out <= 64'b0010011010111000101000111011001010101011101100001010110000000111; end
            14'd11657 : begin out <= 64'b1010100000111010000110101010010010100101101110111001101101010101; end
            14'd11658 : begin out <= 64'b1010101000001011001000011111100010101001111001100010011100110111; end
            14'd11659 : begin out <= 64'b0001101000111011001010110011111110101000011011110010001111101110; end
            14'd11660 : begin out <= 64'b1010100101101010000101110000001110011000101000010010001101111001; end
            14'd11661 : begin out <= 64'b0010101100010011000111001010100010100100011000111010101010011111; end
            14'd11662 : begin out <= 64'b1010011100101110001001100010010010101011010011111010010111111110; end
            14'd11663 : begin out <= 64'b1010101001110000101010101101010010101000000101000010101001110010; end
            14'd11664 : begin out <= 64'b1010101100110001101000110000001000100000001101111010010100001111; end
            14'd11665 : begin out <= 64'b0010000100001000001001101100001100101100000100001010010110011000; end
            14'd11666 : begin out <= 64'b1010101011111000001010010010101110101001001101001010101001101000; end
            14'd11667 : begin out <= 64'b1010100011111011001010000000000100100111010110100010100000100001; end
            14'd11668 : begin out <= 64'b0010000011110000001001010111000010101010100010110010101001111100; end
            14'd11669 : begin out <= 64'b0010000011011111101010000000011000101010000110100001010110011011; end
            14'd11670 : begin out <= 64'b0010100000110110001000001110001110101011110100100001110101001100; end
            14'd11671 : begin out <= 64'b1010100010011110100111100010110010101011101000100010001001101100; end
            14'd11672 : begin out <= 64'b0010000000001000001000111101010010101001001000100010100101101000; end
            14'd11673 : begin out <= 64'b1001111000101010101010101101100100100100000010110010010111010011; end
            14'd11674 : begin out <= 64'b0010011010100101001010100011100110100000100100111010101110011110; end
            14'd11675 : begin out <= 64'b0010101100010011001010100001010000101010110000010010100010000111; end
            14'd11676 : begin out <= 64'b0010101110110010101001010111101100100111011010110010011111101101; end
            14'd11677 : begin out <= 64'b1010100100111010001001000110010010101010000101001010011101011001; end
            14'd11678 : begin out <= 64'b1010100111011100001000110100101100101001001111010010100011010100; end
            14'd11679 : begin out <= 64'b0010100010000111001010000011011010101000011000111010011111010010; end
            14'd11680 : begin out <= 64'b0001111000110101001001000011010010101010111101000010101100010100; end
            14'd11681 : begin out <= 64'b1001110001101001001001101000101110101011010101110010101010010000; end
            14'd11682 : begin out <= 64'b0010100110111111100111011100110110101001000000110010100100000111; end
            14'd11683 : begin out <= 64'b0010000001101100101010000011011100100100100111101010010001010011; end
            14'd11684 : begin out <= 64'b0010101111111010001000000110000100101010111101101010100011010010; end
            14'd11685 : begin out <= 64'b0010101001011000101001000000010000100101101000010010101001111110; end
            14'd11686 : begin out <= 64'b1010000111110001101000110100100110100100110100101010101010001111; end
            14'd11687 : begin out <= 64'b0010100000001111100110001000110000011101010110110010100110111010; end
            14'd11688 : begin out <= 64'b0010010111000001001001010110100010100110100000101010101110101010; end
            14'd11689 : begin out <= 64'b0010100000011010001010110101100110100111111100110001111001001001; end
            14'd11690 : begin out <= 64'b0010000010100000101000110010001100100101111000001010001000010001; end
            14'd11691 : begin out <= 64'b1010011110000100001010001100100010101001100111010010101100111001; end
            14'd11692 : begin out <= 64'b0010011001110010001010001111000110101001101000110010011000001110; end
            14'd11693 : begin out <= 64'b0010010011001110101001111110000000101010000110111001110100001011; end
            14'd11694 : begin out <= 64'b0010001011100101101001100011101100101011110001001010101001011101; end
            14'd11695 : begin out <= 64'b0010001110000011001010010111110110101010100101101010101000010111; end
            14'd11696 : begin out <= 64'b1010101101011000101000001101011000101010011001000010010001101100; end
            14'd11697 : begin out <= 64'b0010010000000100001010100010000010100111101100100010101101111001; end
            14'd11698 : begin out <= 64'b1010000000010110100110100101110000101010111100000010101000000101; end
            14'd11699 : begin out <= 64'b0010100111000000101001000100110110101010110010111010011001111101; end
            14'd11700 : begin out <= 64'b0010100011101110001010110111101100100001011011101010100101101101; end
            14'd11701 : begin out <= 64'b1010101101110011001001011110111100101001111001000010101011110110; end
            14'd11702 : begin out <= 64'b1010100000110110101001111111011000101000100011110010101101011101; end
            14'd11703 : begin out <= 64'b0010100001001000000111010101111010101011100110110010001100011010; end
            14'd11704 : begin out <= 64'b0010101001001010101000100111111110100101100011100010101011111100; end
            14'd11705 : begin out <= 64'b1010010011101110101010010100010000100101010000011010010100011011; end
            14'd11706 : begin out <= 64'b1001101110111101001010011000010010100100101011110010100111001100; end
            14'd11707 : begin out <= 64'b1010011001011000101010010100111010101001010011010001111100011111; end
            14'd11708 : begin out <= 64'b1010101001110100000111010100101110101011101111000001011110101000; end
            14'd11709 : begin out <= 64'b0010100101111110001010001001110110100001101001100001110001000100; end
            14'd11710 : begin out <= 64'b0010100000101000001001001110000010011111000000110010101110101111; end
            14'd11711 : begin out <= 64'b1010101000100011101010100000011110100010111000010010100010011011; end
            14'd11712 : begin out <= 64'b0010101011101001100110011101010100100100000111100010100011000101; end
            14'd11713 : begin out <= 64'b1001011101001011101010100000111010100110100100000001100101111110; end
            14'd11714 : begin out <= 64'b0001111011000100001010100111011010100001110000100010011111110110; end
            14'd11715 : begin out <= 64'b1010001000001111001001111110110100101001001101001010010100100001; end
            14'd11716 : begin out <= 64'b1010101001101010000110110101101010100101101100101010101111001100; end
            14'd11717 : begin out <= 64'b1010100101110001001001010111111000101000111000011010001110011000; end
            14'd11718 : begin out <= 64'b0000110100000000101010011100010100100001011100001010010011100111; end
            14'd11719 : begin out <= 64'b0010101001100001101000111000001110011100010101001010000101000100; end
            14'd11720 : begin out <= 64'b0010010011111111100111100111011100101001011001110010101110111110; end
            14'd11721 : begin out <= 64'b0010101101110000100110000111001110101010100111010001101001010101; end
            14'd11722 : begin out <= 64'b1010011101100001101001101111110000100110101110110010100111001000; end
            14'd11723 : begin out <= 64'b1010010110100101100110000100100110101000111111000010001111111100; end
            14'd11724 : begin out <= 64'b1010011011011100001010000000101010011100100111110010010101101100; end
            14'd11725 : begin out <= 64'b0001010011100000101010011100111110101010000001111010100100000110; end
            14'd11726 : begin out <= 64'b1010001000000110101010110111001110101000000000111010011110111100; end
            14'd11727 : begin out <= 64'b1010010110110010101010001101111010101000010011100010010011001000; end
            14'd11728 : begin out <= 64'b0010010111010010101010111000000100101000111100111010101000010101; end
            14'd11729 : begin out <= 64'b0010011001011100101001010010110000100101010010100010010000011001; end
            14'd11730 : begin out <= 64'b0010101110101100101010101101011010101000111110111010010010111011; end
            14'd11731 : begin out <= 64'b0010001110001101001000001011000110101001111000110001111001010111; end
            14'd11732 : begin out <= 64'b1001110000110011001001110111110000100101010111100010101111100010; end
            14'd11733 : begin out <= 64'b0010011110111011001010011010100110100011111001000010101010101010; end
            14'd11734 : begin out <= 64'b0001101000001101001010000011111110101011100101101001101000110011; end
            14'd11735 : begin out <= 64'b0010100000011111001000011110000010100100010001111010010011000000; end
            14'd11736 : begin out <= 64'b1010011101000001001010010100010010101001100001101010000001001000; end
            14'd11737 : begin out <= 64'b1010011100001000001011000010111000100000110011010010011000100011; end
            14'd11738 : begin out <= 64'b0000110000110100101010100001101100100101010111100010101100000011; end
            14'd11739 : begin out <= 64'b0010101011111100000111100000110110101000000110001010010011100010; end
            14'd11740 : begin out <= 64'b0001111100011101101001001101011100101010010011000010110000010010; end
            14'd11741 : begin out <= 64'b1001110111010001101001101101101100011111011101000001111010101100; end
            14'd11742 : begin out <= 64'b0010101111001101001001000001011000101010110011011010100010001001; end
            14'd11743 : begin out <= 64'b0010100001100100101010000111001010100111110010100010010001000000; end
            14'd11744 : begin out <= 64'b0010101011001011001001011000000000101000010001010010100011011101; end
            14'd11745 : begin out <= 64'b1010000100100100000111001101001010100111110101010010100000000100; end
            14'd11746 : begin out <= 64'b0010101011110010000111010101100110101010010101001010001011000000; end
            14'd11747 : begin out <= 64'b1010100101111101001001000000001100101011011000110010100111101000; end
            14'd11748 : begin out <= 64'b0010100011111100101010000001010110101001011100101010101111001011; end
            14'd11749 : begin out <= 64'b1010011011101110001010111011010010101010000100001010011101000100; end
            14'd11750 : begin out <= 64'b0010101100000110001000100111111110101001011100001010101011000101; end
            14'd11751 : begin out <= 64'b1010101000011001000100011001000000101010100011010010100011101101; end
            14'd11752 : begin out <= 64'b0010011001010010001010011011001110101011010111111010100111001101; end
            14'd11753 : begin out <= 64'b0010010000110010101010000011000100100011110100000010010001100110; end
            14'd11754 : begin out <= 64'b1010100101010001001000101000010000101011010100101010100111100011; end
            14'd11755 : begin out <= 64'b1010011001001001001010000010001100101010001111110000101010100100; end
            14'd11756 : begin out <= 64'b1000111000101100101010110000000100100000100001011010100000101001; end
            14'd11757 : begin out <= 64'b0010001000001010101001101001010010010110100011100010011101100101; end
            14'd11758 : begin out <= 64'b0010010000101100000101100111110000011001010111010010101001001010; end
            14'd11759 : begin out <= 64'b1010100111010001101010011110110010100011000001000010100100101110; end
            14'd11760 : begin out <= 64'b0010100001111011001001110001111100101001000000001010001010110101; end
            14'd11761 : begin out <= 64'b0010101111001111001001001010010000100110011001111010100011100101; end
            14'd11762 : begin out <= 64'b1010001101001111101000101111111000101010110011000010100101010010; end
            14'd11763 : begin out <= 64'b1010100100110100001010001101010110010111100011100010011100101011; end
            14'd11764 : begin out <= 64'b1010101111100101001001110100001000100011100111001010000011011000; end
            14'd11765 : begin out <= 64'b0010000011011111101001000110001000011010100101010010100111000110; end
            14'd11766 : begin out <= 64'b0010011111010010001010111101011010101011001100110010100110001001; end
            14'd11767 : begin out <= 64'b0010100001010010101010111001010000100100001110100010101011011010; end
            14'd11768 : begin out <= 64'b0010010010010011001010111101110100100000001111100010100101010100; end
            14'd11769 : begin out <= 64'b0010011101100000101010100110111010010001101110101010101100001101; end
            14'd11770 : begin out <= 64'b1010001000110001101010001010100000101001001000101001101011000010; end
            14'd11771 : begin out <= 64'b0001111010000100001010010001111000101000100000001010100101001101; end
            14'd11772 : begin out <= 64'b0010010010100100001010100100001010100101110000110010100110101111; end
            14'd11773 : begin out <= 64'b0010101010000011101001111011000010101010000011010010100101101100; end
            14'd11774 : begin out <= 64'b0001010001001000100110111100100000100100101100011010101101011111; end
            14'd11775 : begin out <= 64'b1010011011010101000111010111111110101000101001010010001000100110; end
            14'd11776 : begin out <= 64'b1010100111110011001010000000000110101010100111010010100101001111; end
            14'd11777 : begin out <= 64'b0010000010000010001010011100111000101001001111000010001100000010; end
            14'd11778 : begin out <= 64'b1001010011011100101010101000110110101001101110001010101101101100; end
            14'd11779 : begin out <= 64'b0010011010000001001010001101110110101000000110101010000001001011; end
            14'd11780 : begin out <= 64'b1010100101100010101000100110110000011111111010110010101001110001; end
            14'd11781 : begin out <= 64'b0010011011100000000100100010001000101000101111001010010111010101; end
            14'd11782 : begin out <= 64'b1010100000100111001000010000110110101010110010100010001001110111; end
            14'd11783 : begin out <= 64'b0010101110011101001010000011111000011011000111100001111111100011; end
            14'd11784 : begin out <= 64'b0010011100011110101000010000001100101010011111101010011000001010; end
            14'd11785 : begin out <= 64'b1010101010001000101010010000000110100001101101111010100111001101; end
            14'd11786 : begin out <= 64'b0010101110011010001010000001101110101001010101100010101000101010; end
            14'd11787 : begin out <= 64'b1010010111000001101001011011000100101001010001001010010010010011; end
            14'd11788 : begin out <= 64'b1010100111000010101000111011011000100001111111110010010010010011; end
            14'd11789 : begin out <= 64'b1010101001000111001000001010101100100000000111000010100000100000; end
            14'd11790 : begin out <= 64'b0010001111011010101000000000011000101000100011000001100110111000; end
            14'd11791 : begin out <= 64'b0010011011011000001001101110010100100110000101101010100110001001; end
            14'd11792 : begin out <= 64'b1010101011010001101010110101101010100000001001000010101100101010; end
            14'd11793 : begin out <= 64'b1010010010011100100110001111101000101001011100000010010001100101; end
            14'd11794 : begin out <= 64'b1010101110001011001000111100110110100111100111100010100101110111; end
            14'd11795 : begin out <= 64'b0010011100101100101010111011101100100101110110010010101001101100; end
            14'd11796 : begin out <= 64'b0010100001110111101000100010111000100011011100111010100010001101; end
            14'd11797 : begin out <= 64'b1010010011111000101001011100011100100111100000000010101111111100; end
            14'd11798 : begin out <= 64'b0010010111111001001010001101001010100111001111100010100100100010; end
            14'd11799 : begin out <= 64'b0010000011010011001001010101011110101000011110011010000100100110; end
            14'd11800 : begin out <= 64'b1010010111010000001010101001100000100101111000011010101010100011; end
            14'd11801 : begin out <= 64'b1010010101000001001010100001101110101000001110101010100011101111; end
            14'd11802 : begin out <= 64'b1010100001010111001001100111010010101010000101011010010111101111; end
            14'd11803 : begin out <= 64'b0010100110010101001000110011000010101001010001111001100101001101; end
            14'd11804 : begin out <= 64'b1010100100101111101010101000101110100000011010101010100111110100; end
            14'd11805 : begin out <= 64'b0010100011011100001010100010101100101001000110101010100010010000; end
            14'd11806 : begin out <= 64'b1010100001010101001010000110100010011110100001111010011111101010; end
            14'd11807 : begin out <= 64'b1010010101100101001010101010011110100111000101101010100110111011; end
            14'd11808 : begin out <= 64'b1001001110011000001010111000001010100011001000101010101000101010; end
            14'd11809 : begin out <= 64'b0010101101110001000111011011111100101000001000000010000101001101; end
            14'd11810 : begin out <= 64'b0010000001111011101010010010100100101100010001111010011110011001; end
            14'd11811 : begin out <= 64'b0001010110111011001010010000011000100110111101100010110001010001; end
            14'd11812 : begin out <= 64'b0010011100000000101000111011101010101000110110010010011110000011; end
            14'd11813 : begin out <= 64'b1010101100100010101000100010001110100110010010100001110001100110; end
            14'd11814 : begin out <= 64'b0010101000000010101000101000001010101001101100011010001010110011; end
            14'd11815 : begin out <= 64'b1010100100110101101001011110011000100110100000010010100101001011; end
            14'd11816 : begin out <= 64'b0010001010011000001010001000110000101000011101111001111010101000; end
            14'd11817 : begin out <= 64'b1010101101100101101010001111000010100101110000010010001010110100; end
            14'd11818 : begin out <= 64'b1010010011010101001001111010100100100100110010101010101010001010; end
            14'd11819 : begin out <= 64'b1010011000011101101011000011000100101000100110011010010011000110; end
            14'd11820 : begin out <= 64'b0001110110001000101001101001000010101000101101110010011100110101; end
            14'd11821 : begin out <= 64'b1010100001011111100111111110001010011010000000010010010000011001; end
            14'd11822 : begin out <= 64'b0010010111111000101010010010111110101001010001111010100101110110; end
            14'd11823 : begin out <= 64'b0010110000001111101000101110100000101011001011111001100011010100; end
            14'd11824 : begin out <= 64'b0010011101111101101000100101000000100100010111010010100010000001; end
            14'd11825 : begin out <= 64'b1010101000010100101010011010001000011010100110111010010011111101; end
            14'd11826 : begin out <= 64'b1010100001111100000111011001111100101001110000100010001010010101; end
            14'd11827 : begin out <= 64'b0010100000010000101010000100111110100001110101000010100101001110; end
            14'd11828 : begin out <= 64'b0010001010110010001010000111101010101010110010000010011101011101; end
            14'd11829 : begin out <= 64'b1001100111100010101010000010111000100111000000101010100010001101; end
            14'd11830 : begin out <= 64'b1010010001010110001001100000001110100011001100101010100101111010; end
            14'd11831 : begin out <= 64'b1010100001110110001010000011101010101010100110101001101010110100; end
            14'd11832 : begin out <= 64'b0010001100011001101010100010000100100000110010000010100100110100; end
            14'd11833 : begin out <= 64'b0010100000110101001010111111000110011001011000001010101110001101; end
            14'd11834 : begin out <= 64'b0010010101010101101001111111110110101010010010011010000010001010; end
            14'd11835 : begin out <= 64'b0010100000100111000111010110010010100100001001011010101101111011; end
            14'd11836 : begin out <= 64'b0010101001111010001010100001100000100100110101010010011011100001; end
            14'd11837 : begin out <= 64'b1010010111110011101001111000101010101001011001100001110110011000; end
            14'd11838 : begin out <= 64'b0010100110001101100111000110011110101100000001111010011001010100; end
            14'd11839 : begin out <= 64'b1001101100100110001010000110101110011110011010101010100011100010; end
            14'd11840 : begin out <= 64'b1010010010010111101010010101011100101010111111101010010011101100; end
            14'd11841 : begin out <= 64'b1010101010111110001010111100010000101100001100100001010011110111; end
            14'd11842 : begin out <= 64'b1001101100110001101010000101101110101000110110011010010011110110; end
            14'd11843 : begin out <= 64'b0010101001111011001001100100100010101100010100100010100111101010; end
            14'd11844 : begin out <= 64'b1010100011001000001010010100011010101000110001001010100011111100; end
            14'd11845 : begin out <= 64'b1001110110001101001010111111010110101011100010101010000101001111; end
            14'd11846 : begin out <= 64'b0010100001101011001010010110101110100110101101110010011001001111; end
            14'd11847 : begin out <= 64'b0010000110011000001000001110001010101000100010111010100011001001; end
            14'd11848 : begin out <= 64'b1001111110100101001001011000000110101001111111011010101100100011; end
            14'd11849 : begin out <= 64'b1010000011100010101010010110001100101001110000000010101011000001; end
            14'd11850 : begin out <= 64'b1010011000111110001010101001011100100101100100111010010001111000; end
            14'd11851 : begin out <= 64'b1010101011011111101001101010011000101000001100110010010100000001; end
            14'd11852 : begin out <= 64'b1010100101110001001010010001001100101001001100101010101111101000; end
            14'd11853 : begin out <= 64'b0010101101000110101010011101011110101001101010101010100001111100; end
            14'd11854 : begin out <= 64'b1010011001100100100111101101100000100001111100100010010010111101; end
            14'd11855 : begin out <= 64'b0010000110110100101010110100001010101010110100011010101010010001; end
            14'd11856 : begin out <= 64'b1010011100010011101001110100110000100001010000010010001010011111; end
            14'd11857 : begin out <= 64'b1010000010001111101001111000001110101001011011111010101100011100; end
            14'd11858 : begin out <= 64'b1010100011011000001000001001110000100000011110011010000110110111; end
            14'd11859 : begin out <= 64'b1010100000010101001010110000011000100101001111001010101111010011; end
            14'd11860 : begin out <= 64'b1010100111010110001010001110001100101010000001111010101110100000; end
            14'd11861 : begin out <= 64'b0010000001100101001011000010110010100010011010101010101010111111; end
            14'd11862 : begin out <= 64'b0010101011110000001010111110100010100011101100001010011100010000; end
            14'd11863 : begin out <= 64'b0010100100000000001010111000000010101000101101111001111011110010; end
            14'd11864 : begin out <= 64'b1010010101010110101010110000101100101011001101010010101001101111; end
            14'd11865 : begin out <= 64'b0010001100100010100111011000010010100101010011110010001110111011; end
            14'd11866 : begin out <= 64'b0010011010100001100101010000010100101001001011000010101000101011; end
            14'd11867 : begin out <= 64'b0010101101000011101010110101100010101001000001101010101111111001; end
            14'd11868 : begin out <= 64'b1001110011110011101000011011011000100001100110100010010111001111; end
            14'd11869 : begin out <= 64'b1001000101111100101010010110000110100100011011110010101101100010; end
            14'd11870 : begin out <= 64'b0010011001001111100111110101101110101001011101000010011101100100; end
            14'd11871 : begin out <= 64'b0010010011000001001001010101010000100111001110000010101001101110; end
            14'd11872 : begin out <= 64'b1010001011110101101010011110111110100101111101100010010100111101; end
            14'd11873 : begin out <= 64'b0010100101000000000111101001000100101010100100001010100100100110; end
            14'd11874 : begin out <= 64'b0010011000010011001000100010010000101011011101111010101111000011; end
            14'd11875 : begin out <= 64'b0010000111001100001010011001001010101010101000001010011010111111; end
            14'd11876 : begin out <= 64'b1010101110000111101001100101001100101001110010101010100010110010; end
            14'd11877 : begin out <= 64'b1010100100000001001001001001000100101000110011011010100110100111; end
            14'd11878 : begin out <= 64'b1010011000111111101010000010111110101001011110110010100011000110; end
            14'd11879 : begin out <= 64'b1001010111010111001001000100000100100111111100100010100100001001; end
            14'd11880 : begin out <= 64'b0010101011100110101001111110100110100011110000110010010100110010; end
            14'd11881 : begin out <= 64'b0010011101110111001001010011011010101001000011100010011011101110; end
            14'd11882 : begin out <= 64'b0010001011011101101000110110101010101010110001101010101010111000; end
            14'd11883 : begin out <= 64'b0010011101100101101000110111010100100110100010010010101100100001; end
            14'd11884 : begin out <= 64'b1010101101111110001001101100000010100101010101111010100000111000; end
            14'd11885 : begin out <= 64'b0010010111110010001000110100011110100111101010001001111000100111; end
            14'd11886 : begin out <= 64'b1010100011010110001000000110001110100101011100100010101111000010; end
            14'd11887 : begin out <= 64'b0010001111011110001010111010100110100001001101010010100110111001; end
            14'd11888 : begin out <= 64'b0010001001010000101010010110101000101001111100110010100111111110; end
            14'd11889 : begin out <= 64'b0010100000111000000011100111010110011111000111100010010111000101; end
            14'd11890 : begin out <= 64'b1010010001001001001000001010011110101000010111110001010010001110; end
            14'd11891 : begin out <= 64'b1010101001001011001001001010011110100000010101110010011101110110; end
            14'd11892 : begin out <= 64'b1010001110010110001010110000111010010101011011011010101010001111; end
            14'd11893 : begin out <= 64'b0010101110010011001010000111110010101001110001011010001000011101; end
            14'd11894 : begin out <= 64'b1010000010010010101001100110011010100100101101101010010101010111; end
            14'd11895 : begin out <= 64'b1001111011100000000111001001001010101011000000001010011101110011; end
            14'd11896 : begin out <= 64'b0010101010010000101010111110001000100000001101111010101100100101; end
            14'd11897 : begin out <= 64'b0010011101010100001000000100111100010110010011100010100000000110; end
            14'd11898 : begin out <= 64'b0010101010111000101001011100101010010110010110101010011111001101; end
            14'd11899 : begin out <= 64'b0010010011001000101001001110100110011100101000111010101111000000; end
            14'd11900 : begin out <= 64'b0010010100001111001010110100110100100111010100001010000001000101; end
            14'd11901 : begin out <= 64'b1010100101011010101001010110000110011110001010001010100101010101; end
            14'd11902 : begin out <= 64'b0010100100100110001010001100101000101010110100001010011101000111; end
            14'd11903 : begin out <= 64'b1010001110110111000111010010011010101010101110011010100100000000; end
            14'd11904 : begin out <= 64'b0010010100111110001001100110100100101001000011000010011001100100; end
            14'd11905 : begin out <= 64'b1010101000000001001000101001001100101100010101101010100100000111; end
            14'd11906 : begin out <= 64'b0010001101010010001001110111110010101000101011110001111111000011; end
            14'd11907 : begin out <= 64'b1010010100101100001001100110101010011001110101111010010001000101; end
            14'd11908 : begin out <= 64'b1010100100001110101010111100101010100110110100001010011000101010; end
            14'd11909 : begin out <= 64'b0010001011000110000111110111000100100000100001011010100111011000; end
            14'd11910 : begin out <= 64'b0010101110111110101010000110000100100101011010101010000001101010; end
            14'd11911 : begin out <= 64'b0001111010011001001010110000010110100100101011100010011111010101; end
            14'd11912 : begin out <= 64'b1010010001100010101010011001010110100110001111111010100011011101; end
            14'd11913 : begin out <= 64'b0010101101110010101001110100011110101001101001110010010000000001; end
            14'd11914 : begin out <= 64'b1010100000001000101010101100110000101011010011110010000000101000; end
            14'd11915 : begin out <= 64'b1001011001100001101000100110000100101010100110011001111011011000; end
            14'd11916 : begin out <= 64'b1010101001011000101010001101100000101000001011101010011101101111; end
            14'd11917 : begin out <= 64'b0001101100111011001010101110101110101010110101001010100011000111; end
            14'd11918 : begin out <= 64'b0010001010000110001010000011010010101011111101001010101100100100; end
            14'd11919 : begin out <= 64'b1010010010100100101000100010001000011000001001101010101110111111; end
            14'd11920 : begin out <= 64'b1010010111111001101001110000101010100000100000001010100000011000; end
            14'd11921 : begin out <= 64'b0001111110101111001010001011011010101001001010010010101010101100; end
            14'd11922 : begin out <= 64'b0010100001111101001001010010101100101001000001100010010110101011; end
            14'd11923 : begin out <= 64'b1010110000011000001010000001100100011100001111011010101111001101; end
            14'd11924 : begin out <= 64'b1010101011110101001010100011111100101010110111001010100100101111; end
            14'd11925 : begin out <= 64'b1010000100111011101001101111100110101000111001010010011101001001; end
            14'd11926 : begin out <= 64'b1010000011101111101010100001110000100100100100110000001111101111; end
            14'd11927 : begin out <= 64'b1010000110110101101010111100100100101001111111101010101100010100; end
            14'd11928 : begin out <= 64'b1010011110101010001000001101100110101010010000100010011101001100; end
            14'd11929 : begin out <= 64'b0010101001000111000111001011111010101000011101011010101100111101; end
            14'd11930 : begin out <= 64'b1010100010001110101001010100010110101010100111010010000101110100; end
            14'd11931 : begin out <= 64'b0010100111101010101001011100010000100001100100011010100000000010; end
            14'd11932 : begin out <= 64'b0010010010011100001001111001010110101000000110000010101111110011; end
            14'd11933 : begin out <= 64'b1010011000110111001010100110100010101000010010101010100101010100; end
            14'd11934 : begin out <= 64'b0010100010110011001001000101111100101011010011111010100110001010; end
            14'd11935 : begin out <= 64'b0010101100110100100111011011001000101010111011000010100100111010; end
            14'd11936 : begin out <= 64'b0010000011101011001001000010001110101011111110100010010110001001; end
            14'd11937 : begin out <= 64'b0010000010011101100110110011110000101000011011010010010101000100; end
            14'd11938 : begin out <= 64'b1010101110100001101001101100101010101001101110001010010111001111; end
            14'd11939 : begin out <= 64'b1010010111001011001001010000001100100101000000101010011111100111; end
            14'd11940 : begin out <= 64'b1010101000000001100111100111000110101000110100111001100001001111; end
            14'd11941 : begin out <= 64'b1010101010101100001001011001010110100100101101000001110000111101; end
            14'd11942 : begin out <= 64'b1010011101101010101010000110010110100011110001001010001111101011; end
            14'd11943 : begin out <= 64'b0010100111000100101010001000101100100110010111010010101110011101; end
            14'd11944 : begin out <= 64'b1010100001010000101001011111110110101010011100111010011111100001; end
            14'd11945 : begin out <= 64'b1010100111100001101010001000101110101001001001100010011100100001; end
            14'd11946 : begin out <= 64'b0010101000110011101010000110101010101001101011110010101111001001; end
            14'd11947 : begin out <= 64'b1010010011010001101001000000101010101011100110111010010111001000; end
            14'd11948 : begin out <= 64'b1010101010100000001010010011001000100001000110100010010100100100; end
            14'd11949 : begin out <= 64'b1010011110111100001001000010011100101001110101101010100000100111; end
            14'd11950 : begin out <= 64'b1010101010011000101010010010101110100111110110011010100001001101; end
            14'd11951 : begin out <= 64'b1001110110010010001010110000001100011100101101000001100000111011; end
            14'd11952 : begin out <= 64'b1010101011101000001001011111100100100110110111110010101011111101; end
            14'd11953 : begin out <= 64'b0010100001001100001010001001100110100110111010010010100111111000; end
            14'd11954 : begin out <= 64'b0010010011000101001010101110100110011010111111111010101100001000; end
            14'd11955 : begin out <= 64'b1010100101001101001010011110101110101001010111100010100011001101; end
            14'd11956 : begin out <= 64'b0010100100000011001001011101010110100001010111011010101010010011; end
            14'd11957 : begin out <= 64'b0010100001110010001001011111000010101011000111000010101111110011; end
            14'd11958 : begin out <= 64'b0010101100110100001001110011100110101010111101000010001100001000; end
            14'd11959 : begin out <= 64'b1001111010000110100110011010000000101010100100110010011010011101; end
            14'd11960 : begin out <= 64'b0010101000111100001001101101000100100100010100100001111010010100; end
            14'd11961 : begin out <= 64'b1010101100001111100111011001110110100100010000011010101111100111; end
            14'd11962 : begin out <= 64'b0001011110010011001010000010001010101010100001000010100101011111; end
            14'd11963 : begin out <= 64'b0010101110000001001011000101001010100110100100011010001110110011; end
            14'd11964 : begin out <= 64'b1010011011000001001010111000111000100001000101101010100010010110; end
            14'd11965 : begin out <= 64'b1010101110000100001001110101101010010110001011111010101000000001; end
            14'd11966 : begin out <= 64'b0010000001010110101010111101110110100001011101000010010001101000; end
            14'd11967 : begin out <= 64'b1010010100001101101001111011111000101000100010001010101001001010; end
            14'd11968 : begin out <= 64'b1010101101001000101010001011011100100011010011011010100000100000; end
            14'd11969 : begin out <= 64'b0010101111000111001000000100000100100011001011101010100010000111; end
            14'd11970 : begin out <= 64'b0010011100001101101010011011100010101011111100001010100010100001; end
            14'd11971 : begin out <= 64'b0010101001100001101010100100111000101010001111100010010001000111; end
            14'd11972 : begin out <= 64'b0010100001000010001010011111011000100100001110110010101101001001; end
            14'd11973 : begin out <= 64'b0010100011011101001001000101111000100110011001110010100111111010; end
            14'd11974 : begin out <= 64'b1010101110101011001001001101101000100101011111101010100000101011; end
            14'd11975 : begin out <= 64'b0010010100010000101010001010110010101000000001100001111010011111; end
            14'd11976 : begin out <= 64'b1001101000000010001010110001010100101010110011110010101001010001; end
            14'd11977 : begin out <= 64'b1010010111111100001000000000111110011000001100101010100111011001; end
            14'd11978 : begin out <= 64'b1010100111100100001001001001101000100011100000111010100011101011; end
            14'd11979 : begin out <= 64'b0010010101011010001001010000101000101011001111101010010111010010; end
            14'd11980 : begin out <= 64'b1010101010001111001010001101011000101010111001010010000110011111; end
            14'd11981 : begin out <= 64'b0010001100101110000111111011101110101000011101000010101011000111; end
            14'd11982 : begin out <= 64'b1010100010011110001010011000100000100111001000101010011111000001; end
            14'd11983 : begin out <= 64'b1010100100111001001001000010110000101100001100110010010110111001; end
            14'd11984 : begin out <= 64'b0010100011111110001010001110011110101011110010001010011111101001; end
            14'd11985 : begin out <= 64'b1010011101010101001001101000000000100101111010010010100110111101; end
            14'd11986 : begin out <= 64'b0010010001000011100110100010000010101010001111111010011111001100; end
            14'd11987 : begin out <= 64'b0010101110110111101010111011010010100000010000111010101100011000; end
            14'd11988 : begin out <= 64'b0010000011010100101010000101001100011111001001110010100110100101; end
            14'd11989 : begin out <= 64'b1010011001000101101000100110001010101000110111111010011000011000; end
            14'd11990 : begin out <= 64'b1010011001100110001010011100000010101001110000010010010011001011; end
            14'd11991 : begin out <= 64'b0010010000011110001000011000110000101000111111101010100010010000; end
            14'd11992 : begin out <= 64'b1010000100001000001010001001001000101011110101000010010010001111; end
            14'd11993 : begin out <= 64'b0010000010001010001010011000000110101001011011110010000110101101; end
            14'd11994 : begin out <= 64'b1010100101010111101000010111101110011110111111101010010111101000; end
            14'd11995 : begin out <= 64'b1010100010101111100010100111110010100001101001011010100100101000; end
            14'd11996 : begin out <= 64'b1010101111111001001010011011110000101010000000011010101101000000; end
            14'd11997 : begin out <= 64'b1010101110011101001010111110000010100101011001011001101011010110; end
            14'd11998 : begin out <= 64'b0010101011010001101010111111010010101011000010101001111000101111; end
            14'd11999 : begin out <= 64'b0010000001101001001010010011100100101001111111111010101100001011; end
            14'd12000 : begin out <= 64'b1010011110110111001010101111011010101000000110111010100001101110; end
            14'd12001 : begin out <= 64'b1010010100100101001010010011011010100011001100111010100101000011; end
            14'd12002 : begin out <= 64'b0010000111000000001010100001001100101011100010110010010001010101; end
            14'd12003 : begin out <= 64'b1010010011001011101010101001101000101000011000111010000111010101; end
            14'd12004 : begin out <= 64'b1010100011010100101001011010000100101011010011101001000111011100; end
            14'd12005 : begin out <= 64'b1010101111111101101001000000011010100110010110101010010011000111; end
            14'd12006 : begin out <= 64'b1010100010010110100110010001011010100100011011010010101110110110; end
            14'd12007 : begin out <= 64'b0010100011100010100111000111011110101010000100000010011001011101; end
            14'd12008 : begin out <= 64'b0010100111100000101010100010001100101001000011110010101011100101; end
            14'd12009 : begin out <= 64'b1010100101101011101010101001000000101001000000010010000010100100; end
            14'd12010 : begin out <= 64'b0010000000100100001010001001100100011001010110001010101110010110; end
            14'd12011 : begin out <= 64'b0010011100100011101001100101111110101010001010110001101101111101; end
            14'd12012 : begin out <= 64'b1010101011100001101001101010110100100111001000111010101100111100; end
            14'd12013 : begin out <= 64'b1010100000011001101010001000000000101011000010100010010110011001; end
            14'd12014 : begin out <= 64'b1010101100101110101010001001000010100100011011000010101100110000; end
            14'd12015 : begin out <= 64'b1010010000001100001011000011000010100100100110100010101011000100; end
            14'd12016 : begin out <= 64'b0010100110001011001010011100111000101011000101011010100000111010; end
            14'd12017 : begin out <= 64'b0010101000011101101001100111110010101000000110001010001011100011; end
            14'd12018 : begin out <= 64'b0001111010000110101010000111010010100101000111100010101010000100; end
            14'd12019 : begin out <= 64'b1001110010111100101010010001111100101011100110100010100001011111; end
            14'd12020 : begin out <= 64'b0010011011010010001001010011100110101011110000110000001001011011; end
            14'd12021 : begin out <= 64'b0010100000111010001010011110110000101011101001000010101001111110; end
            14'd12022 : begin out <= 64'b1010011001101111001000100010011110100101111110101010101011100100; end
            14'd12023 : begin out <= 64'b1010101000001110100111101110100110011110111000101001101011101100; end
            14'd12024 : begin out <= 64'b0010100000000000101001010110000110101001100010001010101011100111; end
            14'd12025 : begin out <= 64'b0001101000111011001010100010001010101010010100001010011010101100; end
            14'd12026 : begin out <= 64'b1010101000101110001001000010110010101010011101111010101101101111; end
            14'd12027 : begin out <= 64'b1010010110010000000101010001100110100011111011101010011001100001; end
            14'd12028 : begin out <= 64'b1010010101110100001000100000101110100110011101100010101010001100; end
            14'd12029 : begin out <= 64'b1010001001010001001010010010100100100110010010010001011111001100; end
            14'd12030 : begin out <= 64'b1010101011111100001001100010010110101010100101011010100111011011; end
            14'd12031 : begin out <= 64'b1010000101111000001001000111110100100001110111110010000010001111; end
            14'd12032 : begin out <= 64'b0010101001011011001010100010110010101010110010010010011111100111; end
            14'd12033 : begin out <= 64'b0010101000010010001001011010110010100101010111000010100011111010; end
            14'd12034 : begin out <= 64'b0010101110110001001010111100011110101000101000010001110011100010; end
            14'd12035 : begin out <= 64'b1010000000001011101001011100010100100011110111010010011000010010; end
            14'd12036 : begin out <= 64'b0010000100111010101010011110110010101010100010000001010101100101; end
            14'd12037 : begin out <= 64'b1010100000001000101010111110010000101000111111010010101011111010; end
            14'd12038 : begin out <= 64'b1001110010101010001001101111100010100110111100100010010000000001; end
            14'd12039 : begin out <= 64'b0010101100100101001010011100101010101001011001000010101010010111; end
            14'd12040 : begin out <= 64'b0001100011001111001000110101010100100101010011001010011011011000; end
            14'd12041 : begin out <= 64'b0010101110010011001010000000100100100000100010011010101111010101; end
            14'd12042 : begin out <= 64'b0010001000101110101001001101111100101011100011101010100011111101; end
            14'd12043 : begin out <= 64'b1010010111001000001001101001011000101010111110001010011001001010; end
            14'd12044 : begin out <= 64'b0010100100000101101001110011010110101011011100111010101010101101; end
            14'd12045 : begin out <= 64'b1010100001011111101010010011101010011111111001101010101010001100; end
            14'd12046 : begin out <= 64'b1010001111111000101010011100000110101001110010101010000011110010; end
            14'd12047 : begin out <= 64'b0010011110111110001010100000101100101000001000011010100110101100; end
            14'd12048 : begin out <= 64'b0010011111010001101001000001010010101010110010101010000000001111; end
            14'd12049 : begin out <= 64'b0001000111001000001010100001100110101010000111111010100110110001; end
            14'd12050 : begin out <= 64'b1010010100111111101001110011010100101001001001000010100110010010; end
            14'd12051 : begin out <= 64'b0010001001100001001010011111111100101010100110011010101001110111; end
            14'd12052 : begin out <= 64'b1010101100111001001010101000011100100111110101111010100100110011; end
            14'd12053 : begin out <= 64'b0010011011011010101010100001101110011110001100100010100011000001; end
            14'd12054 : begin out <= 64'b1010001111101001101000001101111110001100111101010010010001000001; end
            14'd12055 : begin out <= 64'b0010101011111000101010110111100110101010001010010010010000001101; end
            14'd12056 : begin out <= 64'b1010101000111101001010101011101110100100001000001010011100101100; end
            14'd12057 : begin out <= 64'b0001101011010110001010100110111010100000101101000001010110011000; end
            14'd12058 : begin out <= 64'b0010101100111010101010000110010010100001111101001010101100000010; end
            14'd12059 : begin out <= 64'b0010010101010001001010110101111000011110110101010010000100111111; end
            14'd12060 : begin out <= 64'b1010100000010000001010110000110010011100100111110010001110001010; end
            14'd12061 : begin out <= 64'b1010000101111101101010101001010100101011001011001010101110111100; end
            14'd12062 : begin out <= 64'b0010010010111010001010001001001000100111100010101001010100010000; end
            14'd12063 : begin out <= 64'b1010101100111100101001010110001100101001001110000001100010100111; end
            14'd12064 : begin out <= 64'b0010010010001100101000000110010010100100010101010001111110010111; end
            14'd12065 : begin out <= 64'b1010000110010101001000111111111100100011010000110010001011101111; end
            14'd12066 : begin out <= 64'b1010100011010001001001000011110110101011110100110010100011111010; end
            14'd12067 : begin out <= 64'b0010101010010101101010111100001100011110100011100010011000010110; end
            14'd12068 : begin out <= 64'b1010010110001101001001001001101010101000001001110010100010010010; end
            14'd12069 : begin out <= 64'b1010101111010011101010111111111010101011100110111010100000010001; end
            14'd12070 : begin out <= 64'b1010101111110000001010110001000110100101111111001010010000011010; end
            14'd12071 : begin out <= 64'b1010100110000100101010011110000100100001010101010010100011000011; end
            14'd12072 : begin out <= 64'b1010100111110010100010000110110010011101001111111010101001110000; end
            14'd12073 : begin out <= 64'b1010010011111101001010101000100010100100111000111010011110100100; end
            14'd12074 : begin out <= 64'b0010101010011100101001010111101100100111101000001010001000111001; end
            14'd12075 : begin out <= 64'b1010101110100110101001101101111010100111010111101010000011010100; end
            14'd12076 : begin out <= 64'b1010100010010100001001101100010010101011110011001010011001101100; end
            14'd12077 : begin out <= 64'b0010010110001001101010010100011110100100100100100010100100101111; end
            14'd12078 : begin out <= 64'b0010100011110011001010010011100000011000001111011010011111111111; end
            14'd12079 : begin out <= 64'b1010000010101000101010000101001110101000110101101010001001000011; end
            14'd12080 : begin out <= 64'b1010100111001110101000100010101100100001110101100010101101010100; end
            14'd12081 : begin out <= 64'b1010001100110111101000000010100010101000000000011001100011010001; end
            14'd12082 : begin out <= 64'b1010101101010110100101000100011000100110111111100010100000110011; end
            14'd12083 : begin out <= 64'b1010110000100101101000111010011100101000111000100010010100011000; end
            14'd12084 : begin out <= 64'b0001111110111000001010000111001000101011000100010010010000011000; end
            14'd12085 : begin out <= 64'b0010101001010000000100001011100110100110001001010001100001000011; end
            14'd12086 : begin out <= 64'b1010100100010100101010011110001100100101111000001010011011011010; end
            14'd12087 : begin out <= 64'b1010011110010011000111110010100010100101111111010010100101010000; end
            14'd12088 : begin out <= 64'b1010000110110000001000100100011010101011111100110001011000101111; end
            14'd12089 : begin out <= 64'b1001010100110000101010110100000000011101110100110010101010000010; end
            14'd12090 : begin out <= 64'b1010010100001101101010111001011010100111011101101001110000011110; end
            14'd12091 : begin out <= 64'b1010100001010000001001001001001010101010010100100010100100011011; end
            14'd12092 : begin out <= 64'b0010011011000001101001111000101110100000100111110010101100001101; end
            14'd12093 : begin out <= 64'b1001110010011111101001111011001000101000001100110010011100111100; end
            14'd12094 : begin out <= 64'b0010101010101110101001101010110000010001000100110010101110101011; end
            14'd12095 : begin out <= 64'b0010000001011100101001010011001100101010000010110010001011000111; end
            14'd12096 : begin out <= 64'b0001100100000011101010001110011110101000101110111010101100100010; end
            14'd12097 : begin out <= 64'b0010001111110001001001000110000000101001110111000010101110011001; end
            14'd12098 : begin out <= 64'b0010000110010011001001110000001110101000010110100010101111010011; end
            14'd12099 : begin out <= 64'b0010010110110011101010001100100010101010110101100010000001111110; end
            14'd12100 : begin out <= 64'b1010101101100101001010111011000100100100000010101010101100111111; end
            14'd12101 : begin out <= 64'b0010101101101010001001010111101000101010010110010010000000101100; end
            14'd12102 : begin out <= 64'b0010101011011010101010011010001000101011111100110010100011110111; end
            14'd12103 : begin out <= 64'b0001110011010100100111001001011000011110001011111010001111101111; end
            14'd12104 : begin out <= 64'b1010101001100001101001111000011000100111111011010010101100110111; end
            14'd12105 : begin out <= 64'b1010100101111101001010111100010110101000001101010010101101011000; end
            14'd12106 : begin out <= 64'b0001001110011011000111110011100010101010110110111001111001010001; end
            14'd12107 : begin out <= 64'b0010101000011100000111111110010100101010110001100010101011110100; end
            14'd12108 : begin out <= 64'b0010100110001011101010110110010100100100111111100010100010011000; end
            14'd12109 : begin out <= 64'b0001100010000011101001100001000010100000011011100010101010011000; end
            14'd12110 : begin out <= 64'b0010001101111111001010111111010100100010110000001010010110111011; end
            14'd12111 : begin out <= 64'b1010010110001000101010010101101000100000000110001010101011011010; end
            14'd12112 : begin out <= 64'b0001111111101111101010110101000110011111100101101010100010001011; end
            14'd12113 : begin out <= 64'b0010000000101000101010011000011000101011000101101010101100011001; end
            14'd12114 : begin out <= 64'b0010100111100100001000111001010100101001011111110001110101110100; end
            14'd12115 : begin out <= 64'b0010100011010101001001111110110110000101100111101010011111100100; end
            14'd12116 : begin out <= 64'b1001100010011011001001011001000000101000101110010010101111101000; end
            14'd12117 : begin out <= 64'b1010101010001110001010011100101100100101101011110010101100100100; end
            14'd12118 : begin out <= 64'b1010101110001000101001110110100110100101111100001010100010011100; end
            14'd12119 : begin out <= 64'b0010000011100110001010110110110000101010000101111001111001110101; end
            14'd12120 : begin out <= 64'b1010100010000100001001100101011100101000110010011010100101011111; end
            14'd12121 : begin out <= 64'b1010000011011101101000111101011010101010110100010010100001101101; end
            14'd12122 : begin out <= 64'b1010100010000110001010000111011100100100001000111010011000000010; end
            14'd12123 : begin out <= 64'b0010011010000100001010100011011000100010110011100010000011000110; end
            14'd12124 : begin out <= 64'b0010101001001111101000010000000000101011011110011010000110110000; end
            14'd12125 : begin out <= 64'b0010100101010111001010100110011100100011001101101010011101110100; end
            14'd12126 : begin out <= 64'b1010100110111010101001011100101100101011010001010010100110001010; end
            14'd12127 : begin out <= 64'b0010011111010001100110100010001110100101100111100010010001010000; end
            14'd12128 : begin out <= 64'b1010100110000111001010100000100010101010000010111010000000010001; end
            14'd12129 : begin out <= 64'b1010100000100001101000101010110010011110001111100010101001111000; end
            14'd12130 : begin out <= 64'b0001110111000110001010000011010000101010101011110010010101001110; end
            14'd12131 : begin out <= 64'b0010001110110001001010010111101000101010001100011010101100011111; end
            14'd12132 : begin out <= 64'b0010011010101111101010001100111100100001000110011010100001111101; end
            14'd12133 : begin out <= 64'b0010000010110010101010001001000100101001010011000010100100011101; end
            14'd12134 : begin out <= 64'b0010011010000001001010110110111110101011100111011001000000110111; end
            14'd12135 : begin out <= 64'b0010011000100101001000100011010010101000110110010010101011000110; end
            14'd12136 : begin out <= 64'b0010011101000101001001110000110110100011110000000010010001010000; end
            14'd12137 : begin out <= 64'b1010101101100101001010011010011000101000000100001010011110101000; end
            14'd12138 : begin out <= 64'b1010010000100111101001001101010000101011011001111001111001011101; end
            14'd12139 : begin out <= 64'b0010010011101001101001110000011010101000001101010010011110011100; end
            14'd12140 : begin out <= 64'b0010101011000110001001111111110010011111011100101001100100100110; end
            14'd12141 : begin out <= 64'b1010011100100000101001000011110000100011101101100001111000011110; end
            14'd12142 : begin out <= 64'b0010101000101010001010111101101100011101000000010010001111111000; end
            14'd12143 : begin out <= 64'b0001110101010001001000011011000110101011000100100010100011101001; end
            14'd12144 : begin out <= 64'b1010101011011101101000101010110000100011101111111010100101111011; end
            14'd12145 : begin out <= 64'b0010010111000111101001000010111010100000101100110010101110111001; end
            14'd12146 : begin out <= 64'b1010101010011111101010010101000100100100001100110010101010100011; end
            14'd12147 : begin out <= 64'b0010101001001011001000111011000000100001010100100010101111111111; end
            14'd12148 : begin out <= 64'b0010101100011110101001100001101100011110100000001010010100110001; end
            14'd12149 : begin out <= 64'b1010100110110000001010000001000100100110010011000010001100110111; end
            14'd12150 : begin out <= 64'b1010101000111101101010100010011110011111011011110010100101000011; end
            14'd12151 : begin out <= 64'b1010011111101110101001010010010010101011011110001010100111100000; end
            14'd12152 : begin out <= 64'b0010101100000000000110000001110110101011001111001010101010011001; end
            14'd12153 : begin out <= 64'b1010011110101000001000100110100010100101101110011010000001001000; end
            14'd12154 : begin out <= 64'b1010100101011110001001101110100000101001101110010010011110111011; end
            14'd12155 : begin out <= 64'b1010100111010101001001010101110000101011100111001010010011100001; end
            14'd12156 : begin out <= 64'b1010100000110001101001001001101000101000010010011010001010001010; end
            14'd12157 : begin out <= 64'b1010100001101101101010000000001100100010010000011001110001001010; end
            14'd12158 : begin out <= 64'b0010001111001001001001101111010110101001010111111010100100100001; end
            14'd12159 : begin out <= 64'b1010101011111110100111110001101110100100111101110010100010101010; end
            14'd12160 : begin out <= 64'b1010101011100101001010010000001000101001010110001010001111101011; end
            14'd12161 : begin out <= 64'b1010100010010101000111111100010100101010010101001010101001000111; end
            14'd12162 : begin out <= 64'b1010001001010000101000000101000100101011111000101010101010000000; end
            14'd12163 : begin out <= 64'b1010010101101001101001011111010000010100110101110010000111100000; end
            14'd12164 : begin out <= 64'b0010101011110110001001111110110100101010010001101010101001110110; end
            14'd12165 : begin out <= 64'b1010100110111101101010000111000010100100111110110010011100011110; end
            14'd12166 : begin out <= 64'b0010101001110100101010001000110110101010111000110010100010010000; end
            14'd12167 : begin out <= 64'b1010001110001001001001011100001010100100101110001010000110010100; end
            14'd12168 : begin out <= 64'b1010101001011001101000110000100110100100001010111010101101000100; end
            14'd12169 : begin out <= 64'b1010100011101110101010100011110000101001101100110010000010100110; end
            14'd12170 : begin out <= 64'b0001100011000010001001011111100010101001101101111010010000001010; end
            14'd12171 : begin out <= 64'b1010100011101010101000111100011000011100001010001010000100110001; end
            14'd12172 : begin out <= 64'b0010011101000110101001111000011110101011011011001010100101110110; end
            14'd12173 : begin out <= 64'b1010101001111000101001010101101000101001111010110010011001111101; end
            14'd12174 : begin out <= 64'b0010100110111010100111101110101110010000000001110010010111111100; end
            14'd12175 : begin out <= 64'b1010000110101000101001010111011110101010101010100010011010011001; end
            14'd12176 : begin out <= 64'b0010100100010001001001010001110100101010101110110010000010111010; end
            14'd12177 : begin out <= 64'b1010100000000111001010110100100110101000110111011010101011110000; end
            14'd12178 : begin out <= 64'b0010101101001010001010100011001100100000101011011001101000111011; end
            14'd12179 : begin out <= 64'b0010011011010110001001100111101010100101100011011010100001000100; end
            14'd12180 : begin out <= 64'b1010101100010010101001110000001100101001111001000010101110010001; end
            14'd12181 : begin out <= 64'b1010100101110100001010011001101010100111010011110010100000011111; end
            14'd12182 : begin out <= 64'b1010100100100100001010011000001010101001101001101010011000100011; end
            14'd12183 : begin out <= 64'b0010011100101001001001011101110100101001110011100010011101011101; end
            14'd12184 : begin out <= 64'b0010101110010000001001101001010000011000001001000010010100100100; end
            14'd12185 : begin out <= 64'b0010101100100111101001010101101100100010101001001010100010011011; end
            14'd12186 : begin out <= 64'b0001100101111111001001110111000000101010111110000010011110101111; end
            14'd12187 : begin out <= 64'b1000110011110111101001110101011110100111101011100010010101111110; end
            14'd12188 : begin out <= 64'b0001110100101000100101010000110000101001010110010010011000001010; end
            14'd12189 : begin out <= 64'b0001110101111011001001110001010110101000000000011010100100101001; end
            14'd12190 : begin out <= 64'b0010001011111011001010101010111110101010111001010010010110011100; end
            14'd12191 : begin out <= 64'b1010011000101101001001110111000110101011110000100001011110100101; end
            14'd12192 : begin out <= 64'b1010010000011110101010010111101010101010011000110010011001110110; end
            14'd12193 : begin out <= 64'b1010010000100101001010110110000110100111100000011010100100101000; end
            14'd12194 : begin out <= 64'b1010011100111101101010000000011000101001101000001010100111010101; end
            14'd12195 : begin out <= 64'b1010000001000011001010000111011010100111110011100010011001001101; end
            14'd12196 : begin out <= 64'b1001111011000001001010011010100000100100110010110010101110000101; end
            14'd12197 : begin out <= 64'b0001010110111011101010100111111100101011111001001010010111001011; end
            14'd12198 : begin out <= 64'b1010000111000000101000100001100010100001110100111010101000001001; end
            14'd12199 : begin out <= 64'b0010011111011110101000000111001100101010000111010010101111111010; end
            14'd12200 : begin out <= 64'b0010000101100101000110010001100110101001110001001010100110100111; end
            14'd12201 : begin out <= 64'b1001101000000011001001000010111110101000000111001010010111001000; end
            14'd12202 : begin out <= 64'b0001011110110011101001110100111010101010000010100010101010001011; end
            14'd12203 : begin out <= 64'b1010100001011001101010100000100110100100100110001010100001001111; end
            14'd12204 : begin out <= 64'b1010100110011001101000000011111010100000100000101010100111010101; end
            14'd12205 : begin out <= 64'b0010001000001000101010001101111010100011001111001010100010100110; end
            14'd12206 : begin out <= 64'b1010011111110110001010101000001000101011110001111010010010001111; end
            14'd12207 : begin out <= 64'b1001000111100010101000101110001100101000110100000010100111001100; end
            14'd12208 : begin out <= 64'b0010110000010001101010100100101000100111111111101010010101111111; end
            14'd12209 : begin out <= 64'b1010010001100110001001110001101000100101100001001010101110010111; end
            14'd12210 : begin out <= 64'b0010100111111000001001110100010000101011001111011010011111101101; end
            14'd12211 : begin out <= 64'b1010101101110100001010111111011010101001001111110010010110011001; end
            14'd12212 : begin out <= 64'b0010010010011010101001011000010000101011001010100010101010010111; end
            14'd12213 : begin out <= 64'b1010101100010010101010101111000000100101001101001010011101101011; end
            14'd12214 : begin out <= 64'b0010100011101011001010111110101110100110110000101010100101001110; end
            14'd12215 : begin out <= 64'b1010100100011101001010010100010010101001011101101010100000100000; end
            14'd12216 : begin out <= 64'b0010010101011000001001111001001100101011111001001010100111010110; end
            14'd12217 : begin out <= 64'b1010000001000101001000011000110110011111000000000010011111110100; end
            14'd12218 : begin out <= 64'b0010101110101110001001100011110110101010100000000010010100001110; end
            14'd12219 : begin out <= 64'b0001100100001100101010100100111000011101111111101010101000010000; end
            14'd12220 : begin out <= 64'b1010101000001000101010100011010010101000100101010010001111010111; end
            14'd12221 : begin out <= 64'b1010101111001010101010111111010000101000010010001010001110111010; end
            14'd12222 : begin out <= 64'b0010100101101011001010011011100110100010001111100001111000101000; end
            14'd12223 : begin out <= 64'b1010100011011000100111000101011100100011001100111010100010010011; end
            14'd12224 : begin out <= 64'b0010100011000111101001000111101110100001011001101010000011111110; end
            14'd12225 : begin out <= 64'b1010011111101100001010101111000100101011111001111010101101110011; end
            14'd12226 : begin out <= 64'b0010100010000011101001101001001010100010011010110001101010111111; end
            14'd12227 : begin out <= 64'b0010011010000110001001000110000010101011010110001010101010000111; end
            14'd12228 : begin out <= 64'b1001101110110011101010100011011000101011001010100010010101100100; end
            14'd12229 : begin out <= 64'b0010100010110110001010011000000010101011101011100010011001111000; end
            14'd12230 : begin out <= 64'b0010000101010110101001101011010100100010100000011010100011100010; end
            14'd12231 : begin out <= 64'b1010100011001111001010011111011100101000000110001010100111010000; end
            14'd12232 : begin out <= 64'b0010101011010010101010000100000100101000011000100010100010110100; end
            14'd12233 : begin out <= 64'b0010100111100100100110001011001100101011010011101010010011111001; end
            14'd12234 : begin out <= 64'b0010101101101001001000110011100110011100000001001010100111001000; end
            14'd12235 : begin out <= 64'b1001111100111001001001100101101110100000011111111010010000001101; end
            14'd12236 : begin out <= 64'b1010100101010000001001000110101000101000010101001001111000010101; end
            14'd12237 : begin out <= 64'b0010100111100000001000111101000010100001111110110010010011100000; end
            14'd12238 : begin out <= 64'b0010011010011110101001100110110100101011100111001010001000100011; end
            14'd12239 : begin out <= 64'b0010101101011011101000111101000010101011011011000010100101101010; end
            14'd12240 : begin out <= 64'b0010100101100001001010000010000100100010101110100001010111111011; end
            14'd12241 : begin out <= 64'b0010011110001101001010000011101000101001011001101010011110011101; end
            14'd12242 : begin out <= 64'b1010011000101110101010101111011100101001100010000010100110110000; end
            14'd12243 : begin out <= 64'b1010101000101111001010000110010010101011110001100010101110110011; end
            14'd12244 : begin out <= 64'b1010010111001111000111010001101010101011001101110010000011100010; end
            14'd12245 : begin out <= 64'b0010101001001110101010010011000100100100110110010010100111101111; end
            14'd12246 : begin out <= 64'b1010010111111101101010001011000100101010101010001010011110111100; end
            14'd12247 : begin out <= 64'b0010101000001010001010100011010110100110001001000010011101000100; end
            14'd12248 : begin out <= 64'b0010101110110000101010100111100100101001111110110010100100010011; end
            14'd12249 : begin out <= 64'b1010010111000011101010101010111010100101000111101010011100000001; end
            14'd12250 : begin out <= 64'b0010100010110011001001111111101000100000001111011010011001111000; end
            14'd12251 : begin out <= 64'b0010101010011111001010111001110010100100010001001010101101110000; end
            14'd12252 : begin out <= 64'b0010101011000110001001010111010010101001111011110010100111100011; end
            14'd12253 : begin out <= 64'b0010101010001111101010001110101000100101110111001010100110101010; end
            14'd12254 : begin out <= 64'b1010010110001101101000110101001110100110010100110010101100110011; end
            14'd12255 : begin out <= 64'b1010110000110010101001001000101100101010100100111010100001000010; end
            14'd12256 : begin out <= 64'b0010001111100110100110000000011110101001101011001010001000010011; end
            14'd12257 : begin out <= 64'b0010110000100101101010001011000010100010101101111010000101000010; end
            14'd12258 : begin out <= 64'b0010001110100000101000000011101100101000011100101010100111110110; end
            14'd12259 : begin out <= 64'b0010100101011110001000010110111110011000011001000001110111010101; end
            14'd12260 : begin out <= 64'b1010010111000010001010001011111010100111000111111010010110001001; end
            14'd12261 : begin out <= 64'b0001100011110100001010101001001110101000000101100000000111010111; end
            14'd12262 : begin out <= 64'b0010011010001010101001011001110100100111110110011010101011011100; end
            14'd12263 : begin out <= 64'b0010110000010111001010100010111010100110010101010010011001010010; end
            14'd12264 : begin out <= 64'b1010011011110000101001000010001000100111010001101010000100100100; end
            14'd12265 : begin out <= 64'b1010101001101111100111100010111000101000111100001010100000100100; end
            14'd12266 : begin out <= 64'b0010101011000011101010111111111100100101111000000010101001111110; end
            14'd12267 : begin out <= 64'b1010100110001110101010010111101000100100001100001010101111000110; end
            14'd12268 : begin out <= 64'b0010101110010000001010101011001110101011101001010000101010010101; end
            14'd12269 : begin out <= 64'b0001111110010010101010001010010100101011100011001010011110101001; end
            14'd12270 : begin out <= 64'b0010100000100000000010010001111100101001110010101010101001001010; end
            14'd12271 : begin out <= 64'b1010011111110111000101000010000010101010001001001001000111011010; end
            14'd12272 : begin out <= 64'b1001111011011011001010000101111010100111010111010010100011001111; end
            14'd12273 : begin out <= 64'b0001111100100011001000001100101010011001011101011010100000001100; end
            14'd12274 : begin out <= 64'b0010101100001010000111110000010110101010001000100010001110100101; end
            14'd12275 : begin out <= 64'b1010100110011011001001101111100010101010010010101010011000011000; end
            14'd12276 : begin out <= 64'b0010100001001110100110100101011110101000000110010001111111100000; end
            14'd12277 : begin out <= 64'b0001110010100100101010101010001100101011101101111001110000010010; end
            14'd12278 : begin out <= 64'b0010011010111011001000010101101010101001000110101010100001101110; end
            14'd12279 : begin out <= 64'b0010000101001010101000011111101110101011001100001010100101111000; end
            14'd12280 : begin out <= 64'b1010101001000111001010000000001100010000101100010010010000001111; end
            14'd12281 : begin out <= 64'b0010011110011000101001110101100100101011100010101001110110000110; end
            14'd12282 : begin out <= 64'b0010001001100100000110011011100010101011011101011010011001100100; end
            14'd12283 : begin out <= 64'b0001110010001010101010000111111010101001110000111010101001001110; end
            14'd12284 : begin out <= 64'b1010010011001010101010000001010110101010011010001010100110000100; end
            14'd12285 : begin out <= 64'b0010011110010101001001100101101000010011001011010001111101110001; end
            14'd12286 : begin out <= 64'b0010101101111110101010010100010010101011110101010010101110010010; end
            14'd12287 : begin out <= 64'b0001100111000001001010010010100000100101001001001010100100110100; end
            14'd12288 : begin out <= 64'b1010011100010100001001110110101110101001100111011010100111111000; end
            14'd12289 : begin out <= 64'b0010100011100011101010011101001010101000001000010010100110010110; end
            14'd12290 : begin out <= 64'b0010100111111010100111000010100000100100000111111010101111001000; end
            14'd12291 : begin out <= 64'b1010010011000011001001110111000000100001111000000010001001101000; end
            14'd12292 : begin out <= 64'b1010101000100000001001100110100110100000001000101010101001000100; end
            14'd12293 : begin out <= 64'b1010000000101011001010100111110000101001001011110001101100011111; end
            14'd12294 : begin out <= 64'b0010010100001111001000001010111110101010001011001010100101000000; end
            14'd12295 : begin out <= 64'b0010100100110101100111010100110100100110011011000010101100110011; end
            14'd12296 : begin out <= 64'b0010100000110110100111111101011000011111100011010010010001100100; end
            14'd12297 : begin out <= 64'b1010011111110001101010000010100010100010000101101010101011100110; end
            14'd12298 : begin out <= 64'b0010101011011001001001110011011110100111100000111001110110111000; end
            14'd12299 : begin out <= 64'b1010101110000101001010011011001100101001000001100010011011011011; end
            14'd12300 : begin out <= 64'b1010011100110011001001011101100010100111111111000010000110010000; end
            14'd12301 : begin out <= 64'b0010101110111011101010100011010110100110111000110010010110100111; end
            14'd12302 : begin out <= 64'b0010100100011000000111100011101110101010111101000010100110010110; end
            14'd12303 : begin out <= 64'b1010100111101011001000101010011010100100000010010010010100001001; end
            14'd12304 : begin out <= 64'b0010100000110100101010101010110010100011110000110010101101000011; end
            14'd12305 : begin out <= 64'b1010011110000111101010100000010100100111001110100010100100000100; end
            14'd12306 : begin out <= 64'b1010011110111001101010010100110110011111100110001010101000100110; end
            14'd12307 : begin out <= 64'b0010100110100011001010000101111110101000111111000010101010101010; end
            14'd12308 : begin out <= 64'b1010100111111111001010100100101000100101111010010001110110010100; end
            14'd12309 : begin out <= 64'b0001111110011001001010111110110000101001011101101010100001010111; end
            14'd12310 : begin out <= 64'b0001010011111111001001001011110110101010001000101010011101011001; end
            14'd12311 : begin out <= 64'b0010101011001111101001110100011000100001001100110010101100001101; end
            14'd12312 : begin out <= 64'b0010101101100011101001100100000010101011110111011010011111010101; end
            14'd12313 : begin out <= 64'b1010001000101000001000010101000110011100010011010010101100101001; end
            14'd12314 : begin out <= 64'b1010100000101110101001010001100100101001101100001010100100110111; end
            14'd12315 : begin out <= 64'b1010101101010100001010110011011110100101010000011010000111100111; end
            14'd12316 : begin out <= 64'b1010000100110111001010011000010000100111010110000010000010100110; end
            14'd12317 : begin out <= 64'b0010100010111110101010001011000000101000111100010001111011011100; end
            14'd12318 : begin out <= 64'b1010011101011010101010110011110000101000000111001010001110001001; end
            14'd12319 : begin out <= 64'b1001111010011110101010010010000000101000001110000010001110100111; end
            14'd12320 : begin out <= 64'b0010100000000101001001100111110010101001101100111010100000100100; end
            14'd12321 : begin out <= 64'b1010100111110100001001000010011000101010011001101010001100010101; end
            14'd12322 : begin out <= 64'b1010101101101101000111001001110010101000101111011001101000111100; end
            14'd12323 : begin out <= 64'b1010100111110000001010100100110010101000111011111010100010111101; end
            14'd12324 : begin out <= 64'b0010011000110111101000101010000110100111100001010010101111101000; end
            14'd12325 : begin out <= 64'b1010100001111001101000111010111100100100000100110010101111000110; end
            14'd12326 : begin out <= 64'b1010100000010110001000101011101110011011011011101010100100001001; end
            14'd12327 : begin out <= 64'b0010010110011110000110111100000000101000010101010001111100111000; end
            14'd12328 : begin out <= 64'b1010001011111011001010011111001010101000000100011010101001001110; end
            14'd12329 : begin out <= 64'b1010000100101010100111100110111100100110110100111010100000010101; end
            14'd12330 : begin out <= 64'b0010100101110100101010010011110010101001010001110001111010101101; end
            14'd12331 : begin out <= 64'b0010101010000011101000110101001010101011001011001010000010011011; end
            14'd12332 : begin out <= 64'b0010011001100011001000010000011000100111110100110010010110100111; end
            14'd12333 : begin out <= 64'b0010100110100011101010010010111100101011001010011010010000101111; end
            14'd12334 : begin out <= 64'b1010101001110011101000101110100000100111001110001010101101100000; end
            14'd12335 : begin out <= 64'b1010100000111110101010111110110110100000001000010010010111100111; end
            14'd12336 : begin out <= 64'b1010100000011101001001111000100110101001101100100010101001001010; end
            14'd12337 : begin out <= 64'b1010100110100111001010001000111000101011011110001010101110010110; end
            14'd12338 : begin out <= 64'b0010100111011000001001010010111100101001000001110010100100010001; end
            14'd12339 : begin out <= 64'b0010001101000000101010100101100100100000100011100010101100100010; end
            14'd12340 : begin out <= 64'b1010101001001110001000110011010100010101001001110010100101001001; end
            14'd12341 : begin out <= 64'b1010101110000001100111110010000000101001010000011010010101011011; end
            14'd12342 : begin out <= 64'b0001111000110110001010011101010010101011111011101010101101000011; end
            14'd12343 : begin out <= 64'b0001110110000100101010001011010100100101000000001001100101010011; end
            14'd12344 : begin out <= 64'b0010000000110100001001100001101110101000100001001010100010011110; end
            14'd12345 : begin out <= 64'b1010100010101111101001101001110100100110110100001010010001111101; end
            14'd12346 : begin out <= 64'b0001101100001000001000010100011000101011110111010010101000000001; end
            14'd12347 : begin out <= 64'b1010100101111001101010101101100000100100110100111001100010100110; end
            14'd12348 : begin out <= 64'b1010000101111001001000101011010000101010111100101001110001111111; end
            14'd12349 : begin out <= 64'b0010100010111010100101100100000010101010000001101010100000101000; end
            14'd12350 : begin out <= 64'b1010100000101101101001101011010100100100111100011010010011010100; end
            14'd12351 : begin out <= 64'b1001101000010001101010100011000010011101101110111010010010101100; end
            14'd12352 : begin out <= 64'b1010100110110101101001101100011110101010000011000010010101000010; end
            14'd12353 : begin out <= 64'b1010011100110010101001110001111100101001010001011010011100010010; end
            14'd12354 : begin out <= 64'b1010101001000100101001001011101110100110111100111010010101101110; end
            14'd12355 : begin out <= 64'b1010010110111101101000100100010110101010010001000010011001100101; end
            14'd12356 : begin out <= 64'b1010100000100011001010000010111110101010010010001010100100010010; end
            14'd12357 : begin out <= 64'b0010100110101110001010111101000000101001010011011010101100011010; end
            14'd12358 : begin out <= 64'b0010011101011011101001011101001100101000010110101010101011100011; end
            14'd12359 : begin out <= 64'b1010100101000111001001101011010000101001011101001010001100100001; end
            14'd12360 : begin out <= 64'b1010011101010011100110011000111100001001000100000010101111111111; end
            14'd12361 : begin out <= 64'b1010011010011001101010011110000010010100111100010010100101111101; end
            14'd12362 : begin out <= 64'b0010101001011111100101000011011010101001001110000010101100101010; end
            14'd12363 : begin out <= 64'b1010101110010010001010010010110110101011010001000010010011100000; end
            14'd12364 : begin out <= 64'b1010101011010100001001011100000000101010011011101010100001111001; end
            14'd12365 : begin out <= 64'b0010101001100000001010000000001110011011100010101001111101011111; end
            14'd12366 : begin out <= 64'b1010110000001001001010110100110110101010101000110010010011110000; end
            14'd12367 : begin out <= 64'b0010010110010010101000100000001010100010101111100010010011000001; end
            14'd12368 : begin out <= 64'b1010101010110000001010101100100100100101111000001010110000010000; end
            14'd12369 : begin out <= 64'b1010010100001101101010111110101100011110101011010010000111110110; end
            14'd12370 : begin out <= 64'b1010010000101000101000010000000110101001100000100010101000000111; end
            14'd12371 : begin out <= 64'b1010001101100010001010001101111000101010011000101010100000101110; end
            14'd12372 : begin out <= 64'b0010010000000011000101000111000110101011001101110010100100111011; end
            14'd12373 : begin out <= 64'b1010010001000101001001110101000010100100111110101010101010001000; end
            14'd12374 : begin out <= 64'b0001011001011101101001101111100000011000110000011010100010111001; end
            14'd12375 : begin out <= 64'b0010100101000000101010111011001110101000100000100010101101001011; end
            14'd12376 : begin out <= 64'b1010101011000111101010100000001110101011110000011010100011110000; end
            14'd12377 : begin out <= 64'b0010101101000110101001111111111000101001011110110001110001111000; end
            14'd12378 : begin out <= 64'b1010010011011011001001000011010010100111000101011001100001101101; end
            14'd12379 : begin out <= 64'b0001100010110010001001001011000100100111000010000010100001100000; end
            14'd12380 : begin out <= 64'b0010011101100000001000110101101110100111101001000010100100001101; end
            14'd12381 : begin out <= 64'b0010000000101101001001001100100100100100010100011010101011110011; end
            14'd12382 : begin out <= 64'b0010101110010101001000001100100100100001000110110010101010111011; end
            14'd12383 : begin out <= 64'b1010101011000010000111110010110100101000100001010010100010100100; end
            14'd12384 : begin out <= 64'b1010100100101010101010001001000100101000110011111010011000010001; end
            14'd12385 : begin out <= 64'b0010000100111110001001011101111110100100110101001010101001111110; end
            14'd12386 : begin out <= 64'b0010011111101001101001000110111110101000000010011010100101100001; end
            14'd12387 : begin out <= 64'b1010100101111101101010001010110010101000010000101001101011000111; end
            14'd12388 : begin out <= 64'b0010100101101110101000110011111000100010000011100001110000110111; end
            14'd12389 : begin out <= 64'b1010100101101111001010101000000100100011101111111010100110100010; end
            14'd12390 : begin out <= 64'b1010011011001001101010000110001110011000010100110010010100110001; end
            14'd12391 : begin out <= 64'b0001101000111011001010101101111100100110011000100010100001110011; end
            14'd12392 : begin out <= 64'b0010101100001100001010011011000010101001010100111010000000001000; end
            14'd12393 : begin out <= 64'b0010000111001101101010101001000000101000011010110001111001010111; end
            14'd12394 : begin out <= 64'b1010101101001111100000111000000000101000001010000010100010101100; end
            14'd12395 : begin out <= 64'b0010001101010101000110111011001110100110101110000010100011000101; end
            14'd12396 : begin out <= 64'b0010101011010001001010101100101000101001110011000010010100010100; end
            14'd12397 : begin out <= 64'b0010011010100111001001010111001110100000101001110010011101101100; end
            14'd12398 : begin out <= 64'b1010100011111111101010100011001010100010000100110010010100001010; end
            14'd12399 : begin out <= 64'b0010000100010100101001101110011110101001101110101010100010001001; end
            14'd12400 : begin out <= 64'b1010101110010010101010010011110010101001011100010010100101110010; end
            14'd12401 : begin out <= 64'b0010101010011100101010110001100000100101001001101010101110111100; end
            14'd12402 : begin out <= 64'b1010100110111011101010011110110110101011110111000010001010011010; end
            14'd12403 : begin out <= 64'b0010101100000100001010111111010100100110101010001001111001001100; end
            14'd12404 : begin out <= 64'b0010100011010110101010001110010000100110001010001010101000000110; end
            14'd12405 : begin out <= 64'b1010101101010001101010010011011100011111000010110010011110001011; end
            14'd12406 : begin out <= 64'b0010100101000010000111111001100000011110010001011010101110111001; end
            14'd12407 : begin out <= 64'b1010100011100000001001111101111000011010100001110001100010100001; end
            14'd12408 : begin out <= 64'b0010011011000100101010100110011100100100101101101010100001000001; end
            14'd12409 : begin out <= 64'b1001110001110101001010001101100100100000101001010010100110000100; end
            14'd12410 : begin out <= 64'b1010011001001111100101100100110110100101001111100010000100101010; end
            14'd12411 : begin out <= 64'b0010100100100001001010000111101110101011100111101010100110100001; end
            14'd12412 : begin out <= 64'b1010100101100101001010011111000010011110011100000010101100011101; end
            14'd12413 : begin out <= 64'b1010101010000110100110101110011100100100111001101001101101010110; end
            14'd12414 : begin out <= 64'b1010100100101100001010011011110010100101000100101010100010100000; end
            14'd12415 : begin out <= 64'b1010101011101100001001101010111100101010011110000000111111000010; end
            14'd12416 : begin out <= 64'b1010101000010101001000101100111100101010101111100010001111000010; end
            14'd12417 : begin out <= 64'b0010101111100010101010111100100110101011110110100010100010011001; end
            14'd12418 : begin out <= 64'b0010101000101110000111000110110110100110011100110010101000111010; end
            14'd12419 : begin out <= 64'b0010101101111001001010110001100110100111011100100010000111101010; end
            14'd12420 : begin out <= 64'b0010100110100000001010010001100110101001001011111010011000100111; end
            14'd12421 : begin out <= 64'b1010001100011000101001000110010000101000111000001010001101000110; end
            14'd12422 : begin out <= 64'b1010100111110010101001100011011000100101110100010001110000100001; end
            14'd12423 : begin out <= 64'b0001110111101111001010101011100110100111111110000001011001000011; end
            14'd12424 : begin out <= 64'b1010101011010001000110000110010100100111110111100010100111011010; end
            14'd12425 : begin out <= 64'b1010100110011001101010111010101000101010110111000010011000111010; end
            14'd12426 : begin out <= 64'b1001110000101011001000011000000100101001001010101010010010001101; end
            14'd12427 : begin out <= 64'b0010011101110001101010000110101100101011011010110010011000010100; end
            14'd12428 : begin out <= 64'b1010101011011110001010111101011010101000011011001010001101101100; end
            14'd12429 : begin out <= 64'b1010100110011101001010000000011110100110011001001010100100101011; end
            14'd12430 : begin out <= 64'b1010001100111010001010101101010000100011101111110010101000001000; end
            14'd12431 : begin out <= 64'b0001110101110000101000110000000100101010001011011010100100001001; end
            14'd12432 : begin out <= 64'b0010001100001010101001000111011000101001111110100010010000010001; end
            14'd12433 : begin out <= 64'b0010000000001011101010010100100100101010000110010001110000001111; end
            14'd12434 : begin out <= 64'b0010000011011110001010111110011010010101001000111010101111010000; end
            14'd12435 : begin out <= 64'b1001101111100000001010100110101100100111011100001010011111010110; end
            14'd12436 : begin out <= 64'b1010100100001000001001111010110110101011100101110010100100101010; end
            14'd12437 : begin out <= 64'b1010101000010001001010110000000000101010110100000010100011100010; end
            14'd12438 : begin out <= 64'b1010101100010001101010011110000110100101110111111010100110111001; end
            14'd12439 : begin out <= 64'b0010101011010010001010011011101000100010000100000010011011111001; end
            14'd12440 : begin out <= 64'b1001111000001100101001100001100000011000001011011010100100111000; end
            14'd12441 : begin out <= 64'b0010100111011001101001110011100000101000000000101010101010000110; end
            14'd12442 : begin out <= 64'b0010100000110110001000001011001100010011010011100010101010111010; end
            14'd12443 : begin out <= 64'b0010101001101100001010110010010100100111000010101010101101110001; end
            14'd12444 : begin out <= 64'b1010100110100101001010110100001110100100010011111010101011010011; end
            14'd12445 : begin out <= 64'b0001111000011101101001000100111110101001010000101010010000000111; end
            14'd12446 : begin out <= 64'b0010100100101011001010101101000000101001100111100010001100101010; end
            14'd12447 : begin out <= 64'b1010101100010110101010000100100000100010001000000010000010111011; end
            14'd12448 : begin out <= 64'b1010100100010001001010110001100100101010110110011010100100011111; end
            14'd12449 : begin out <= 64'b0010101000101010001010100000011010101000111001111010000001101100; end
            14'd12450 : begin out <= 64'b1001010011001001101001010101000100011111000000010010100011001110; end
            14'd12451 : begin out <= 64'b1010010010111111001010001110101110011100011110010010100000100010; end
            14'd12452 : begin out <= 64'b1010101001111011001001100101001110010111111001001010101111100000; end
            14'd12453 : begin out <= 64'b1001111111110110001010010001111000101001000100011010100010001100; end
            14'd12454 : begin out <= 64'b1001110111100010101010110001001100011000111110010010010100000111; end
            14'd12455 : begin out <= 64'b1010001110111111100110111000110000100101000100001010001011111111; end
            14'd12456 : begin out <= 64'b0010100011010101001010110000100110100110100101111010101110101110; end
            14'd12457 : begin out <= 64'b1010010010101100001010111101100110101011000000000010101110101010; end
            14'd12458 : begin out <= 64'b0010011000110000001010100101111100001110000000011010100010111001; end
            14'd12459 : begin out <= 64'b0010000000110000000110110111001110101010111110110010100011101111; end
            14'd12460 : begin out <= 64'b1010100101110010001010111101011100101000000000010010010100100100; end
            14'd12461 : begin out <= 64'b1010101010100101101010101000000100011111110000110010010101001000; end
            14'd12462 : begin out <= 64'b1010101001000101101001100011111100101011100010111010000100011010; end
            14'd12463 : begin out <= 64'b0010100111001011001010000110111100101000011010111010011100010111; end
            14'd12464 : begin out <= 64'b0010010011111101001010011010101010101001111011011010100011010101; end
            14'd12465 : begin out <= 64'b1010000000111110001010100000011100101001110000101010100110100000; end
            14'd12466 : begin out <= 64'b1010010100111111101010101000111000100101110001001010011100000000; end
            14'd12467 : begin out <= 64'b0010101010101001001001000110011110101001000000110010010001101100; end
            14'd12468 : begin out <= 64'b1010000110010101001010110011001000100100101111100010011011110000; end
            14'd12469 : begin out <= 64'b0001100101011010001010111111110000100101111101110010100001010000; end
            14'd12470 : begin out <= 64'b0010001110000001001000011001110010100111110101101010011011111100; end
            14'd12471 : begin out <= 64'b1010101001000111001010100110100010100010111101111001101000111111; end
            14'd12472 : begin out <= 64'b0010100001111100100111101101010100101001110000000010101000111101; end
            14'd12473 : begin out <= 64'b1010101000110110001010010001110100100001100011110010100010001001; end
            14'd12474 : begin out <= 64'b1010101011110100001010111010000000100101101001011010010111001010; end
            14'd12475 : begin out <= 64'b1001100011111001101010111001001000101011010101011001111011111101; end
            14'd12476 : begin out <= 64'b1010101000010000101000110011011110101001000100101010100110100110; end
            14'd12477 : begin out <= 64'b0010011001110111101001010011100100101001001111001010000100010000; end
            14'd12478 : begin out <= 64'b1001110011110000001001000011110100101010101100010010001010011110; end
            14'd12479 : begin out <= 64'b1010011110101001100010010101100100100101101011010010100100001101; end
            14'd12480 : begin out <= 64'b0010101001101001101010000000000010011101000100101010010110000010; end
            14'd12481 : begin out <= 64'b1010100111100010101010000001110100101000111001101001010110101000; end
            14'd12482 : begin out <= 64'b1010100100111110000111011100000000101010100110110010100111100011; end
            14'd12483 : begin out <= 64'b1010100000001100101001011011111000101011101100100010100111010111; end
            14'd12484 : begin out <= 64'b0001111010101110001010011111110110100100011000100010101110111000; end
            14'd12485 : begin out <= 64'b0001110110011101101000110111011110011110110100100001101111010111; end
            14'd12486 : begin out <= 64'b0001110111011010101001111010001100101010100011100010101101001010; end
            14'd12487 : begin out <= 64'b1010011101100111101000110011110110100101101001110010100010010110; end
            14'd12488 : begin out <= 64'b0010000111110111101010001000010000100111100101101010100110001010; end
            14'd12489 : begin out <= 64'b0010100110101010101001100110011000100111010000000010000001001011; end
            14'd12490 : begin out <= 64'b1010011000011001001010000000111100100100001111111010000001010010; end
            14'd12491 : begin out <= 64'b0010001011110011101001110100100110100010100101110010101000111010; end
            14'd12492 : begin out <= 64'b0001011110010010100111000001111100101010010001100010011010111111; end
            14'd12493 : begin out <= 64'b1010101100011110001010100001001100011101100010110010001111100000; end
            14'd12494 : begin out <= 64'b0010000000011110001010011101000100101010110001011010001010101000; end
            14'd12495 : begin out <= 64'b0001001111001110101010101001010110100010101010011010101111010010; end
            14'd12496 : begin out <= 64'b0001100000110010001010101101110100100000101010111001110001111000; end
            14'd12497 : begin out <= 64'b0010011010100110001001010101110100011100011011010010101110000100; end
            14'd12498 : begin out <= 64'b0010000010000111001010100101101010101011110111010010100010001001; end
            14'd12499 : begin out <= 64'b1010011000011111100011011000000000011101001000000010100011010100; end
            14'd12500 : begin out <= 64'b1010010010101110000110100001110000101010100001101001101100010011; end
            14'd12501 : begin out <= 64'b1010011001000100000111111110001010101010010110110010011100010000; end
            14'd12502 : begin out <= 64'b0010100000111110100110010110111000100110000001100010101100111101; end
            14'd12503 : begin out <= 64'b1001110111001011001001011010011010100110010000100010100100110011; end
            14'd12504 : begin out <= 64'b0010000111010100101001010011100110100100101000101010100000011001; end
            14'd12505 : begin out <= 64'b1010010110000010001010111000110100100100101110100010000110100100; end
            14'd12506 : begin out <= 64'b0010011111011101101010001011010110101001011011001010010001110111; end
            14'd12507 : begin out <= 64'b1010011011100011101010111010101010100100000101001010100100100101; end
            14'd12508 : begin out <= 64'b0010100101101111001010011111011000101010010000110010101111100101; end
            14'd12509 : begin out <= 64'b1010101010000011101001000000000100100101010000110010011010100100; end
            14'd12510 : begin out <= 64'b1001010110001000101001101110110000101010011111111010010000110000; end
            14'd12511 : begin out <= 64'b0010100011001000101000110011111100100010110011110010010010001000; end
            14'd12512 : begin out <= 64'b0010100010010011001001100111100110101010001011010001110011100100; end
            14'd12513 : begin out <= 64'b0010000100111110001000001000001010101001010111110010011101111011; end
            14'd12514 : begin out <= 64'b1010101111001110101010100001001110101010110000101010101010001010; end
            14'd12515 : begin out <= 64'b1010011001111000100111110001101000011101110111101010101101110110; end
            14'd12516 : begin out <= 64'b0010101001010010101000011001011010011101000011001010011111001011; end
            14'd12517 : begin out <= 64'b0010000001100010101001011000101010100001011010000010101010011101; end
            14'd12518 : begin out <= 64'b0010010110000100001001000110100110100101011110000010100111010011; end
            14'd12519 : begin out <= 64'b0010011110010101001000011011110100100111100011100010100101001010; end
            14'd12520 : begin out <= 64'b1001111100000001001001001000001110101010011101100001010000111001; end
            14'd12521 : begin out <= 64'b0010101001001100101010111011111010101010000010011010010010010000; end
            14'd12522 : begin out <= 64'b0010010101000101101010100001101010100101011101101010011010010110; end
            14'd12523 : begin out <= 64'b0010110000001011001010011000000110101001111011101010100100101000; end
            14'd12524 : begin out <= 64'b1010100110111101001000110000011100100111000000100010100001010001; end
            14'd12525 : begin out <= 64'b1010100000100010001010111100000000011000010110110010100011101010; end
            14'd12526 : begin out <= 64'b1010100000011110101000110100000000101000010011110001010100101110; end
            14'd12527 : begin out <= 64'b0001100001001111001000001101010010100010000110110010101100011010; end
            14'd12528 : begin out <= 64'b1010010001101110101000001101110110101011000001001010010110111101; end
            14'd12529 : begin out <= 64'b0010011011100111000110101110001000101010011100101010101011011101; end
            14'd12530 : begin out <= 64'b1010100010101000001010110100011110101000100100001010101111001111; end
            14'd12531 : begin out <= 64'b1010010111011100101010000001111100100111100111110010001111110001; end
            14'd12532 : begin out <= 64'b1010011110100000101010110001101000100100101110111010011110011011; end
            14'd12533 : begin out <= 64'b1001100011111110001010000111110010101001001011000010011010101011; end
            14'd12534 : begin out <= 64'b0010001110010100001010101001101100101011000111101010010111111100; end
            14'd12535 : begin out <= 64'b0010100110011110101010001101010000101011001011001010001100000111; end
            14'd12536 : begin out <= 64'b1001100100001100101001101000100100100111011101110010101110001101; end
            14'd12537 : begin out <= 64'b1010000010111110001001100111111010101001100000110010011001100011; end
            14'd12538 : begin out <= 64'b1010010101010000000111110000011100011111010111110010011011010111; end
            14'd12539 : begin out <= 64'b0010101101011100001010010010101010101001010100110010101010001110; end
            14'd12540 : begin out <= 64'b0010100000111111001001000100010010100111001110000001001000010000; end
            14'd12541 : begin out <= 64'b1001010001010010001001100100001100101010000111011010100100011100; end
            14'd12542 : begin out <= 64'b0010101011001011001010000011101000101001011111100010010111110110; end
            14'd12543 : begin out <= 64'b1010100001100000101001101100110010100100101001110010110000001101; end
            14'd12544 : begin out <= 64'b1010011111110011101001100001101110100010011010111001111111010110; end
            14'd12545 : begin out <= 64'b1010010001001101001010011001111110100110011101001010101110010011; end
            14'd12546 : begin out <= 64'b1010001010001001001010000101101110011101010001000010101111101111; end
            14'd12547 : begin out <= 64'b1010001000010101001001101000001100100110100101010010100010100101; end
            14'd12548 : begin out <= 64'b1010010101101110101001110101000100101010001010100010100111110101; end
            14'd12549 : begin out <= 64'b1010100101010111101010000011011100101011001110111010010101001010; end
            14'd12550 : begin out <= 64'b1010001000001101001010001110001110101010110011000010100001000101; end
            14'd12551 : begin out <= 64'b0010101000000100101010011100100100101000111111011010001100110000; end
            14'd12552 : begin out <= 64'b0010100100000100100110001010100000101000101011010010100101110001; end
            14'd12553 : begin out <= 64'b1010100111001100101001011000001000101000100001110001111101001011; end
            14'd12554 : begin out <= 64'b1010010010001011101011000000000100100110011101011010100001110010; end
            14'd12555 : begin out <= 64'b1001101011110110101001000100000010011110001011010001011000110100; end
            14'd12556 : begin out <= 64'b1010100110100101101010011100111010101000110010100010101011011000; end
            14'd12557 : begin out <= 64'b0001100000110101101010111100110100100011100110001010100111110011; end
            14'd12558 : begin out <= 64'b1010101011010001001010101101100010101000000011100010100010110000; end
            14'd12559 : begin out <= 64'b1010101000000001101010111101000010011010101011111001010111010100; end
            14'd12560 : begin out <= 64'b0010010100100001001010001001001100101000101010101010011101100111; end
            14'd12561 : begin out <= 64'b1010011100001111101001001110000000100011100101111010100001011011; end
            14'd12562 : begin out <= 64'b1010000101011010101001100110010110100101001000100010101110011011; end
            14'd12563 : begin out <= 64'b0001110011001001101001011101101000101010100100000010100111101100; end
            14'd12564 : begin out <= 64'b1010100100011000001010000100010110000011000001001000100110111001; end
            14'd12565 : begin out <= 64'b0010011111000100101001110010101110101100001111011001001000111110; end
            14'd12566 : begin out <= 64'b1001100000110011001010011101011110101010110011011010010011010010; end
            14'd12567 : begin out <= 64'b0010110000011011100011010101001100101001011111001010101111111100; end
            14'd12568 : begin out <= 64'b0010011011011001101010110010110000100100110001101010100011101010; end
            14'd12569 : begin out <= 64'b0010100000100010101010101100111000011110100100010010101010100011; end
            14'd12570 : begin out <= 64'b0010100000100111101010001001111010100011111000011010100010010100; end
            14'd12571 : begin out <= 64'b0001000011101010001010011010011000011001001111111010011000010010; end
            14'd12572 : begin out <= 64'b1010101001101101101010010110000010100111011100100010100111100010; end
            14'd12573 : begin out <= 64'b1010100000110111101000111111000000100000010000110010101110010100; end
            14'd12574 : begin out <= 64'b1010101000101011101001000101010000101011100000000010101111010110; end
            14'd12575 : begin out <= 64'b1001101000100001001001100001110000101010000010111010000111001011; end
            14'd12576 : begin out <= 64'b0010101101111001001000000000110000011001001101100010001010110000; end
            14'd12577 : begin out <= 64'b0010010000000001100110000101001010100110110000010010010100100101; end
            14'd12578 : begin out <= 64'b0010100100001010101001100000011100100010010110011010100110110101; end
            14'd12579 : begin out <= 64'b0010001011101000101010001011101010011011011000101010010000001011; end
            14'd12580 : begin out <= 64'b0010100110100011101010000010111110100100111100100010011010110010; end
            14'd12581 : begin out <= 64'b1010011110111110101010100000000010101011011110100010100000110100; end
            14'd12582 : begin out <= 64'b1010001000111010000111111010110010011001010001010010100000101011; end
            14'd12583 : begin out <= 64'b0001111111110110101010010110111110100010011111111001111100010111; end
            14'd12584 : begin out <= 64'b0010101111001101001001010000100110100001011101011010100010110110; end
            14'd12585 : begin out <= 64'b0010100010001100101000001010101110100110101001110010101110011001; end
            14'd12586 : begin out <= 64'b1010010111010100001001111110110100100010000110011010100000101111; end
            14'd12587 : begin out <= 64'b0010011010011011001010101101100110011110100011100010100101010001; end
            14'd12588 : begin out <= 64'b0010100010110011001010110111100010011101101111001010101000101011; end
            14'd12589 : begin out <= 64'b1001111101110011100101111110101000101010100001011010000001011100; end
            14'd12590 : begin out <= 64'b0010010100111010001010001100101010101010000101100001010100010111; end
            14'd12591 : begin out <= 64'b1010000110000010101001010101010010100101001010011010011110010001; end
            14'd12592 : begin out <= 64'b0010101100010101001010101111010000101000111000110010001010111001; end
            14'd12593 : begin out <= 64'b1010101101111101001010001100100010100100001101110010010100101010; end
            14'd12594 : begin out <= 64'b0010100001101110001001101000111000101000101100101010001100001100; end
            14'd12595 : begin out <= 64'b1010101011110101001010011010101010100100101001001010101011111110; end
            14'd12596 : begin out <= 64'b0010011101010111001001010000011010100111001011111010101111110000; end
            14'd12597 : begin out <= 64'b1010100101000011001010110100101100101010011001101010010010011111; end
            14'd12598 : begin out <= 64'b0010100100011110000110101011101000101001010000001010011111100100; end
            14'd12599 : begin out <= 64'b0001111100110111101010101101000000101010101001010001111110111011; end
            14'd12600 : begin out <= 64'b1010000100011011101010100000001010100010100000010010100110000010; end
            14'd12601 : begin out <= 64'b1010101100110110001010000110001100101010100001111010100100001110; end
            14'd12602 : begin out <= 64'b1010101010000011001001000101110010011101111100011001111111110001; end
            14'd12603 : begin out <= 64'b1010001100111011001000011000010110100110011001001010000110001000; end
            14'd12604 : begin out <= 64'b1010101110010011001010011101011000100110000101110010101000111000; end
            14'd12605 : begin out <= 64'b1010101111000100001010101010011100101000111000000010101010111111; end
            14'd12606 : begin out <= 64'b0010000001100001001010110100110100100101111001001001111000001111; end
            14'd12607 : begin out <= 64'b0010010010111010000110010011001010100000101111100010011100010110; end
            14'd12608 : begin out <= 64'b1010100010011110001010011101011100101011010111011010001001000110; end
            14'd12609 : begin out <= 64'b0010101101010000001010110011011000001100010010111010101011101100; end
            14'd12610 : begin out <= 64'b0010010101010001101000101111010010100110100110110010011101100010; end
            14'd12611 : begin out <= 64'b1010010001001010100110110111100100101001101100111010100000010011; end
            14'd12612 : begin out <= 64'b1010101101001110001010011101000010101001101111100010000000100011; end
            14'd12613 : begin out <= 64'b1001111010011101001000011011000110011111101010011001110101010001; end
            14'd12614 : begin out <= 64'b1010001011001110100111111110011110011010000010100010101101110010; end
            14'd12615 : begin out <= 64'b1010001001100001101010001001000000100110100101000010001001011010; end
            14'd12616 : begin out <= 64'b0010010100011001101010000100111100101010100110110010100101010101; end
            14'd12617 : begin out <= 64'b1010100000110111001001010010110010101011011100000010010110100110; end
            14'd12618 : begin out <= 64'b1001111011111010001001110100101110010001101101100010101111111011; end
            14'd12619 : begin out <= 64'b1010101110011001101010110011101100101011110010011010101011100101; end
            14'd12620 : begin out <= 64'b0010101000010000101001011010010010100100110110010010001111010100; end
            14'd12621 : begin out <= 64'b0010100111101101100100110101100010011110010100011010101100011010; end
            14'd12622 : begin out <= 64'b1010000101101100101001001000110010100011111110101010101101110001; end
            14'd12623 : begin out <= 64'b1001110011101101001010111000101010101000001000100010011011110011; end
            14'd12624 : begin out <= 64'b0010101001101110001010011011010100101010110100110010100011000001; end
            14'd12625 : begin out <= 64'b1010101111000000101001100011010000101000000110111010101011110001; end
            14'd12626 : begin out <= 64'b1010101110010000101010010111101110100000100101111010100110100110; end
            14'd12627 : begin out <= 64'b0010101101111000101010100100111000011001001001001010011111000111; end
            14'd12628 : begin out <= 64'b0001000111010010101010001110100010101000011100110001100100111011; end
            14'd12629 : begin out <= 64'b0010100111101000001010011110101010100100001110101010100011001101; end
            14'd12630 : begin out <= 64'b1010101001100000101001110110100110101000000010100010101000000011; end
            14'd12631 : begin out <= 64'b0010100011011001001010100011011010100011011011100010101011110000; end
            14'd12632 : begin out <= 64'b0010101110011010100111011011111010100110000001010010101100011111; end
            14'd12633 : begin out <= 64'b0010101001011010101010111101110010101010100100011010010011101011; end
            14'd12634 : begin out <= 64'b0010101100100011001000011100010010101011010101100010010001011011; end
            14'd12635 : begin out <= 64'b0010001110110001101010010010001010100010111100101010001100110100; end
            14'd12636 : begin out <= 64'b0010100011000000101010011101110100100111001101011010101001100001; end
            14'd12637 : begin out <= 64'b1001110111001110001010001001101010100101100001001010101101001110; end
            14'd12638 : begin out <= 64'b0001110100100011101010111100001100100100010001001010101100011001; end
            14'd12639 : begin out <= 64'b1010101100010010001001000110110100101010101011000010011010111100; end
            14'd12640 : begin out <= 64'b0010010101100111101001011100111010100110100000101010100000100111; end
            14'd12641 : begin out <= 64'b1010101001101110001000111001010000101011100100111010100010100110; end
            14'd12642 : begin out <= 64'b1010100100000001101010011110000100100110100011001010101010000000; end
            14'd12643 : begin out <= 64'b1010001011100001100111110010000110100011100010001010010001000000; end
            14'd12644 : begin out <= 64'b1010011001110011101010011111101010100110100000111010101001110001; end
            14'd12645 : begin out <= 64'b1010001110111001101001000111110000100101101101000010000000000000; end
            14'd12646 : begin out <= 64'b0010101000000100001001110000110100101011011110001010001101111000; end
            14'd12647 : begin out <= 64'b0010011001000100101000001100010010101010111100010010100011101010; end
            14'd12648 : begin out <= 64'b0010100011101001101010110010111000010100001101100010100111100111; end
            14'd12649 : begin out <= 64'b1010010010110010001010101010001010101011001001101010011010011011; end
            14'd12650 : begin out <= 64'b0010011000010000100111010000001000100100110100001010100100011000; end
            14'd12651 : begin out <= 64'b0001101010011010101001101100110010101010100101111010101011101100; end
            14'd12652 : begin out <= 64'b0010011101011000000111010011010000101010110001011010010010010010; end
            14'd12653 : begin out <= 64'b1010011000010000001010000010101010100000101101000010011100000010; end
            14'd12654 : begin out <= 64'b0010010010111010101010110111111000101010111100100010101010011001; end
            14'd12655 : begin out <= 64'b1010100110100110101010111010001000100110111001111010101000110101; end
            14'd12656 : begin out <= 64'b1010011010100001101001101110110000100100110011110001111101101100; end
            14'd12657 : begin out <= 64'b1010100011000011001010010001000110100011010011111010101001010100; end
            14'd12658 : begin out <= 64'b0010011000100101101010111010001100100001101101000010011101010111; end
            14'd12659 : begin out <= 64'b0010101000101111101010111100000100100110100000010010101010110001; end
            14'd12660 : begin out <= 64'b1010010100100100101001010011110100101000110010101010101010110001; end
            14'd12661 : begin out <= 64'b0010100010011001001001000110100010100011111100101010001011000000; end
            14'd12662 : begin out <= 64'b0010101100011100101010111101100010100101101011111010001001100100; end
            14'd12663 : begin out <= 64'b1010101100000110101000110110010010101000100110000001110101101101; end
            14'd12664 : begin out <= 64'b1010010010100011100111111110000000011101100001111010100100001101; end
            14'd12665 : begin out <= 64'b0010000100001100001010000101001110100111110011001010101110100010; end
            14'd12666 : begin out <= 64'b1001110001011000001010000001100000011111001000100010100000100011; end
            14'd12667 : begin out <= 64'b1010100001100101001010000000001110101010110100011010100100100101; end
            14'd12668 : begin out <= 64'b1010000111001001001000001101110100101001101010000010100010001010; end
            14'd12669 : begin out <= 64'b1010101100100101001010100000100010101000100110101010000111101011; end
            14'd12670 : begin out <= 64'b0010010011001011000110100110110000100000111110111010101000110110; end
            14'd12671 : begin out <= 64'b0010001000111000101001001011001010101001111101001010100010010101; end
            14'd12672 : begin out <= 64'b1010001100001010001010101010011100101000001110000010100010110110; end
            14'd12673 : begin out <= 64'b0010001010000111000111011000101110101001100100110010101011011110; end
            14'd12674 : begin out <= 64'b0010100110101110101000101000001110011101111010110010101000100100; end
            14'd12675 : begin out <= 64'b0010110001010011001010111010001100100111011010101001110000100011; end
            14'd12676 : begin out <= 64'b0010100001000101001001100111001000101000101011000010101001100111; end
            14'd12677 : begin out <= 64'b1010101010100010101000100100010110011111001011111001110101101011; end
            14'd12678 : begin out <= 64'b0010100111000010001010010000001100101010101010110010101010100100; end
            14'd12679 : begin out <= 64'b1010101110011011001010010101000110101011101000010010011111110110; end
            14'd12680 : begin out <= 64'b0010101110011000001010011100101100100111110101010010101001010110; end
            14'd12681 : begin out <= 64'b1010010110001111001001100101001100101000111000000001101010100110; end
            14'd12682 : begin out <= 64'b0001111011100101001001110110011100101010000001100010100011011110; end
            14'd12683 : begin out <= 64'b0010101100101010101010000011001110101000001100101010100000101001; end
            14'd12684 : begin out <= 64'b1010100010101011000111101101000000101000001000110010001101010110; end
            14'd12685 : begin out <= 64'b1010010110001000101001111110100110100101011101011010101101000101; end
            14'd12686 : begin out <= 64'b0010101000001101001010101010101000101000110100110010101110110101; end
            14'd12687 : begin out <= 64'b0010010110100000101010001100000010100100101111010001110001100110; end
            14'd12688 : begin out <= 64'b0010011100001101001001111110101010100000011000100010000000010001; end
            14'd12689 : begin out <= 64'b0010010011101101000111110000010110100111010000011010100100010110; end
            14'd12690 : begin out <= 64'b0010100101111110101010011101000010101011111111101010100010011001; end
            14'd12691 : begin out <= 64'b1000111010011110101001100110000100101010100001101001110010100000; end
            14'd12692 : begin out <= 64'b0010001101001011101001100010100100100100100111100010100000110001; end
            14'd12693 : begin out <= 64'b1010100111111000101010000111110110100110100110100001111100001010; end
            14'd12694 : begin out <= 64'b0010100110101011001010111101111100101000011100110010101100000011; end
            14'd12695 : begin out <= 64'b0010000110110100001001101100000000101010010110110010010001100000; end
            14'd12696 : begin out <= 64'b1010100000000011001001100001110100101000010110010010101110010101; end
            14'd12697 : begin out <= 64'b0010100110011101101010111100111000101011010010001001111011101110; end
            14'd12698 : begin out <= 64'b1010101110101111101001010100010000101011101100001010011000101010; end
            14'd12699 : begin out <= 64'b0010100011001111001010101101111110100100100111100010011001010111; end
            14'd12700 : begin out <= 64'b0010011011001111001010100010010000100100011101010010010100111001; end
            14'd12701 : begin out <= 64'b0010011110101101101010110000011010100101011111010001111001100000; end
            14'd12702 : begin out <= 64'b0010100010100110000111010110100000100110001111000010010011011000; end
            14'd12703 : begin out <= 64'b1010100010100100101001100111011110101010000100110010100100001110; end
            14'd12704 : begin out <= 64'b0010100111110000101010000110010110101011001000101001111010110110; end
            14'd12705 : begin out <= 64'b1000110001010001101000000110011100101000010000000010100101101101; end
            14'd12706 : begin out <= 64'b0010100101101011001010001110011100100101101000111010100101101101; end
            14'd12707 : begin out <= 64'b0010100000100010101010100010110010101010110011000010011111001101; end
            14'd12708 : begin out <= 64'b0010011001000100001010100001111100101011011110010001001010101000; end
            14'd12709 : begin out <= 64'b1010001001001111001001111100111000101011010000101010101100111101; end
            14'd12710 : begin out <= 64'b1010101101111001001010001111111110100111011011110010011100111111; end
            14'd12711 : begin out <= 64'b1010101001110010101001001010011010101100000110101010101001110111; end
            14'd12712 : begin out <= 64'b0010100111111001101001001001001100101000111101101010000111000101; end
            14'd12713 : begin out <= 64'b0010011001111011101001001110011110011110010011011010001111011110; end
            14'd12714 : begin out <= 64'b0010011010001110000111111100100110101011011011110010100111001101; end
            14'd12715 : begin out <= 64'b0010010110000100100100000011111110100001000010100010101011011101; end
            14'd12716 : begin out <= 64'b1001101011101011100111000001111110101010101101000010011000100101; end
            14'd12717 : begin out <= 64'b0010011110010110001010100001001110101010011001000010101011111101; end
            14'd12718 : begin out <= 64'b1010010111100100001010110100100100101000010000111001111011000010; end
            14'd12719 : begin out <= 64'b1010011101010101001010111001010000101001111110000010100111011010; end
            14'd12720 : begin out <= 64'b1010010110111010101001101001111100100110100001011010000010101101; end
            14'd12721 : begin out <= 64'b0010100011100100101010000010000110101010001010111010101101001100; end
            14'd12722 : begin out <= 64'b0010011111000001101010000111110110101000101001101010011110101001; end
            14'd12723 : begin out <= 64'b1010101010001100001010010110100000100100001111111010100100110101; end
            14'd12724 : begin out <= 64'b1010100101001111001010000111110000101010011010100010100101000100; end
            14'd12725 : begin out <= 64'b1010101111000100101010110110011110101100000010101010011100101010; end
            14'd12726 : begin out <= 64'b1001111110100010101010100111011010100111001100011010011010101100; end
            14'd12727 : begin out <= 64'b0010100010000010101010010101011010101001000101000010001111100011; end
            14'd12728 : begin out <= 64'b1010100100001100101010111000011010101010100000101010101111101100; end
            14'd12729 : begin out <= 64'b1010010011010111101001001110001010101000110110000010101001111001; end
            14'd12730 : begin out <= 64'b1010001110111010001010000010000110101100000100010010011100000101; end
            14'd12731 : begin out <= 64'b0010010111011000001010101010000100101100000010100010000011110011; end
            14'd12732 : begin out <= 64'b0010101111011101101001000010010100101000100001101010100100110110; end
            14'd12733 : begin out <= 64'b0001110011101010101010001010011110100000111010010010100001101111; end
            14'd12734 : begin out <= 64'b1010100101010000101010001100011110011001111110010001110010100001; end
            14'd12735 : begin out <= 64'b1010010101101110101001010010010100100100110100101001111110001101; end
            14'd12736 : begin out <= 64'b1010101001110100101001011110010000100011011110100010100000000001; end
            14'd12737 : begin out <= 64'b0010100010100001001001110100100000100111100111011001101110010110; end
            14'd12738 : begin out <= 64'b0010101010110000101010000011000010100010110001111010101000001000; end
            14'd12739 : begin out <= 64'b0010100010011100001001010001100010100100100111010010100001100010; end
            14'd12740 : begin out <= 64'b1001111111000001001010100011000110100001101001001010101001111111; end
            14'd12741 : begin out <= 64'b0010000101000010101000101100101110100100000111010010011111111111; end
            14'd12742 : begin out <= 64'b1010110000110000101000110101010010101001000010100010011101100100; end
            14'd12743 : begin out <= 64'b0010101101011111100110111011000110101010110000010001100100110011; end
            14'd12744 : begin out <= 64'b0010100001101101001010110011111010101010000000001010010010010111; end
            14'd12745 : begin out <= 64'b0010101101000011101010101110000110101001100100101010101001110011; end
            14'd12746 : begin out <= 64'b0010100010111011001000100110011010101011010111100010011100100000; end
            14'd12747 : begin out <= 64'b1010010101001110000110111010111010100110011011100010101100111111; end
            14'd12748 : begin out <= 64'b0001101100110011001001110010100010100111010010001010100110101111; end
            14'd12749 : begin out <= 64'b0010100100111110100111101011111110011100111100100010100101101110; end
            14'd12750 : begin out <= 64'b0010000011100011100111111110101110101001000111100010100100000110; end
            14'd12751 : begin out <= 64'b1010011100101011000111110010110000101001000111000001111010001010; end
            14'd12752 : begin out <= 64'b1010100111000000001010110001100000101011010101011010001110111000; end
            14'd12753 : begin out <= 64'b1010000101010011001010111110010110100101101101011010010100101110; end
            14'd12754 : begin out <= 64'b0010100000001110001010010101001110101000011010010010100110000100; end
            14'd12755 : begin out <= 64'b1010100010101001001001000101010010101010001110010010101010010111; end
            14'd12756 : begin out <= 64'b0010101010110011001010101110000000101011001001000001111011110001; end
            14'd12757 : begin out <= 64'b1001101001111010001010011000001010010000001011010010100010001110; end
            14'd12758 : begin out <= 64'b1010100001011011101001000111111110101001100111000010100011101100; end
            14'd12759 : begin out <= 64'b0010011000101001100111010110100110101001000011100010101011011001; end
            14'd12760 : begin out <= 64'b1001110110101111001001100001111110101011000011000010011000100001; end
            14'd12761 : begin out <= 64'b1010011101100111101000100100000100101011011001101010100000100001; end
            14'd12762 : begin out <= 64'b0010001011100100101010101011110100100000100000000010001111101101; end
            14'd12763 : begin out <= 64'b0010100100111110001001001101010110011110111101110010011000111000; end
            14'd12764 : begin out <= 64'b0001111101100010101010011011000100101011010100100010010111011001; end
            14'd12765 : begin out <= 64'b1010100111110101000100100001101100101000111001101010010111001011; end
            14'd12766 : begin out <= 64'b1010100010011001101010000011111110100010110100000010100010000000; end
            14'd12767 : begin out <= 64'b0010101000000101001000100001010010101011000010000010100110100011; end
            14'd12768 : begin out <= 64'b0010100000110001001001100100001100011101101010100010101111101001; end
            14'd12769 : begin out <= 64'b0010001110000011101001111000010100100001110101000010001000000001; end
            14'd12770 : begin out <= 64'b1010101111001011001001001100011010101001101111011001101010001101; end
            14'd12771 : begin out <= 64'b1010100100001010001010111001001010100001110000110010101001010011; end
            14'd12772 : begin out <= 64'b1010101101101110001010010011001010101000101110100010101010010111; end
            14'd12773 : begin out <= 64'b0010100010011001101010111100100110101001010111010010100001100101; end
            14'd12774 : begin out <= 64'b0010011011111010001000000111110000100001010000101010010011001111; end
            14'd12775 : begin out <= 64'b1010100111001111001001001010010100100111010101100010001001000011; end
            14'd12776 : begin out <= 64'b1010011101111000001011000001001010101000100001110001000101101111; end
            14'd12777 : begin out <= 64'b0010100010111101001000110101100110101010111100100010011101000010; end
            14'd12778 : begin out <= 64'b1001100101111111001000010100011110101010010001101010010101011101; end
            14'd12779 : begin out <= 64'b0010100110001101001010100001110100011001101111011010001010000000; end
            14'd12780 : begin out <= 64'b0010100001000001101000101110011010001001010101001010010010101011; end
            14'd12781 : begin out <= 64'b1010011110111010001000111101011010100101010101101010100101000101; end
            14'd12782 : begin out <= 64'b1010010011110011101010100100000010101001101101010010100101000001; end
            14'd12783 : begin out <= 64'b1010101000101000101010010001001110101000000100000010100110110111; end
            14'd12784 : begin out <= 64'b0010100101010110001010010001000110101001101101110010100011100111; end
            14'd12785 : begin out <= 64'b0010100110101011001010110110010010011110010010111010100000101010; end
            14'd12786 : begin out <= 64'b0010100110100011001000010101111100101010011101010010100000001101; end
            14'd12787 : begin out <= 64'b1010001010000011001010110011110110101010011000110010100011110101; end
            14'd12788 : begin out <= 64'b0010100011010011001001000011010010101001111010011010101010011101; end
            14'd12789 : begin out <= 64'b0010011001001101101010000101001100011100111110011010101101111110; end
            14'd12790 : begin out <= 64'b0010001011010100101001010011011100101010101011110001110110100111; end
            14'd12791 : begin out <= 64'b1010010011011100100110000111000000011010011111000001111100011101; end
            14'd12792 : begin out <= 64'b0010100110100110101001100101101000101011011000100010101010111001; end
            14'd12793 : begin out <= 64'b0010010011000000001010011110011100101011111011110010100000101111; end
            14'd12794 : begin out <= 64'b0010101010110110101001000000000110100010011001000010010111001111; end
            14'd12795 : begin out <= 64'b1010100100111100101000011010001100101000110110100001110011001000; end
            14'd12796 : begin out <= 64'b0010100011111110000110000101101100101000111101011010100010100100; end
            14'd12797 : begin out <= 64'b0010101011101100101001100101100010101001010111000010010011011100; end
            14'd12798 : begin out <= 64'b1010100011111100101000101110110100011100001110101001010011111010; end
            14'd12799 : begin out <= 64'b0010010000010010001001011011001010101011010000110010100101111110; end
            14'd12800 : begin out <= 64'b0010001100111110000111100110110110011111100000110010010100111001; end
            14'd12801 : begin out <= 64'b0010000011001111001011000000001010011010111111111010100101011110; end
            14'd12802 : begin out <= 64'b1010001000100100100010100011101010101010110010011010011000000110; end
            14'd12803 : begin out <= 64'b1010001011001010001001110010000100101100010001001010100101011100; end
            14'd12804 : begin out <= 64'b1010000011001101101000110011010100101000000101101010101101111000; end
            14'd12805 : begin out <= 64'b0010001011101010101001000100000000101001010100001001111011101100; end
            14'd12806 : begin out <= 64'b0010011000100011101010010101110010101010101101111010010110011100; end
            14'd12807 : begin out <= 64'b1010101001001000000111000000111000101011001010111010000111001110; end
            14'd12808 : begin out <= 64'b1010100001001010001010111111010000100010011000000010101110000011; end
            14'd12809 : begin out <= 64'b1010100111111100001010100100111000011111001000110010100011011011; end
            14'd12810 : begin out <= 64'b0010001101001111001000010001101010101000111010010010001110010011; end
            14'd12811 : begin out <= 64'b0010000000110010001010001100101100100100110101100010101010110000; end
            14'd12812 : begin out <= 64'b0010101010000100101010100010010110101001000001011010101010110010; end
            14'd12813 : begin out <= 64'b1010100010011110001010000100101100100001100110011001100110011111; end
            14'd12814 : begin out <= 64'b0010101011100111100111010011111000011110011111010010011111110001; end
            14'd12815 : begin out <= 64'b0010011010000100001010010011101110100110000101110010101011011001; end
            14'd12816 : begin out <= 64'b0010010000101101001001111101001110101010010110101010100000010111; end
            14'd12817 : begin out <= 64'b0010100110001001101010010101111010101100000111101010100000001110; end
            14'd12818 : begin out <= 64'b1010001000110010101011000000101000101010101001011010101011000110; end
            14'd12819 : begin out <= 64'b1010010100100101001001101111111100101001111110100010011000100001; end
            14'd12820 : begin out <= 64'b1010100100101111001010110100011000100101010010001010101010101010; end
            14'd12821 : begin out <= 64'b0010101011011000101001000011100110101011000110010010000111000110; end
            14'd12822 : begin out <= 64'b1010100100011111100111101101100110100100011101110010011111110001; end
            14'd12823 : begin out <= 64'b1010011100101110101010110111001000101011110001100010101111000100; end
            14'd12824 : begin out <= 64'b1010101101000000001001001101010000101010101101011010010010011101; end
            14'd12825 : begin out <= 64'b1010101000000110100111010001110010100101001000111010010101011100; end
            14'd12826 : begin out <= 64'b1010010101110011101010110110001110101010011001001001110010101000; end
            14'd12827 : begin out <= 64'b1010101010010111001010011110101100100100101110000010010011010100; end
            14'd12828 : begin out <= 64'b0010100111011100101010001001011000101000001001100010101001111110; end
            14'd12829 : begin out <= 64'b0010100111001100001010001011110010101010100100001010011100011000; end
            14'd12830 : begin out <= 64'b1010100110101100101010011100011010100101110101110010100010110110; end
            14'd12831 : begin out <= 64'b1010101010111011100111100111111110101001001101000001001101101010; end
            14'd12832 : begin out <= 64'b0010000100000101101010001010001000101001101000101010010110011010; end
            14'd12833 : begin out <= 64'b1010010001100000001001000011100100101011000101000010010001010011; end
            14'd12834 : begin out <= 64'b0010100110101011001001001110001010100000111111011010101011000000; end
            14'd12835 : begin out <= 64'b1010000100001010001000111000101100101010100100010010001100001110; end
            14'd12836 : begin out <= 64'b1010101110000110101010001010111010100101111011111010101100101000; end
            14'd12837 : begin out <= 64'b0010010111110110101000011100011100101011100111110010101000010100; end
            14'd12838 : begin out <= 64'b0010011011001000000110010010001010100111111100110010011010110110; end
            14'd12839 : begin out <= 64'b0010001001001011001010110000010010101010111110001010000000000000; end
            14'd12840 : begin out <= 64'b0010101011111101001001001100011110100010010001000010101011000010; end
            14'd12841 : begin out <= 64'b0010101000101101001010100110111110101000111110011010010001001111; end
            14'd12842 : begin out <= 64'b0010100111110111101010101010110010101010110100011010101010000110; end
            14'd12843 : begin out <= 64'b1010011001101111001001010011000110101001100001111010101000100111; end
            14'd12844 : begin out <= 64'b0010001001001001001010101001000100101011011011101010011100000011; end
            14'd12845 : begin out <= 64'b0010011111110111101010110001101010100100011001000010010101111101; end
            14'd12846 : begin out <= 64'b0010101011010010001010101001011000100110100010000010100001001011; end
            14'd12847 : begin out <= 64'b1010010000001111001010010110111000101011111100010010010101100110; end
            14'd12848 : begin out <= 64'b0010101000010101101010101110111000101011101010001010101111011000; end
            14'd12849 : begin out <= 64'b0010101111001110101001001001110100101010110101101010011110110000; end
            14'd12850 : begin out <= 64'b0010010011110001001001111001000110100111110110101010011001001111; end
            14'd12851 : begin out <= 64'b0001110111111101001000100011011110100101111011010010001101110000; end
            14'd12852 : begin out <= 64'b0010100111001001000110101100010000101010101010011010010010111010; end
            14'd12853 : begin out <= 64'b1001011000111111101010111010011010011000001101001010101101010101; end
            14'd12854 : begin out <= 64'b1010110000001110101010111001010100100110011000011010101010011001; end
            14'd12855 : begin out <= 64'b1010100100000101001010110111010110101010010100101010000001100110; end
            14'd12856 : begin out <= 64'b0010100101011010101010010000101000101001000011010010010111110000; end
            14'd12857 : begin out <= 64'b1001111100001110001010110100010100101001000100001010100101101011; end
            14'd12858 : begin out <= 64'b1010100010010110001001011111100010101010010000010010100101001011; end
            14'd12859 : begin out <= 64'b1001011010011111101010001011010000100010011010000010100101001100; end
            14'd12860 : begin out <= 64'b1010000011111100101001010000100110101100001101011010100110101011; end
            14'd12861 : begin out <= 64'b1010010110011001101010111111110110100101100010010010100010000000; end
            14'd12862 : begin out <= 64'b0010101011000110101010011010000000101011101110001010100010110001; end
            14'd12863 : begin out <= 64'b0010101000010010001001100110110100101001001010010010010101100100; end
            14'd12864 : begin out <= 64'b1010010101110000101010001101001100101011011001011010100000011010; end
            14'd12865 : begin out <= 64'b1010001111101100101010011011011110011100100011110010100011001101; end
            14'd12866 : begin out <= 64'b1010000010001001001010011110110010010010100101110010011111011000; end
            14'd12867 : begin out <= 64'b1010011001110011001001110101010110101011000111000010101010001010; end
            14'd12868 : begin out <= 64'b1010101111110010101010000110100000101000111101000010100110001100; end
            14'd12869 : begin out <= 64'b1010010100101100101010100110001000000000001000001010101101011111; end
            14'd12870 : begin out <= 64'b1010100111000010101001111100111000101010101100111010011001111011; end
            14'd12871 : begin out <= 64'b1010011001000101001001010110110110101010110101100010000101000111; end
            14'd12872 : begin out <= 64'b1010100001001000001001000011010000100100000111111010100010110101; end
            14'd12873 : begin out <= 64'b0010010101110001100110011001100100100100110100010010100000101000; end
            14'd12874 : begin out <= 64'b0010011101001010001001010011100010100110110100110010000111100110; end
            14'd12875 : begin out <= 64'b0010010100100011101000011001000000101011000111110010100001000101; end
            14'd12876 : begin out <= 64'b0010100000101010001001101111111010011110011110011010010011100101; end
            14'd12877 : begin out <= 64'b1001100100001110001010010100110010100100010100001010000001010111; end
            14'd12878 : begin out <= 64'b0010101010010101101001001000010010101000111110011010011111011100; end
            14'd12879 : begin out <= 64'b1010010011101000001001010001110110010110010000000010100110100001; end
            14'd12880 : begin out <= 64'b0010011101101100001000011101101110101001001001101010101111001001; end
            14'd12881 : begin out <= 64'b0010100010001010101001010111001110100011101101000001111110000011; end
            14'd12882 : begin out <= 64'b0010010000100011001001010000110000101010001000111010100111101011; end
            14'd12883 : begin out <= 64'b0010101100111001001010100110001100100001010110000010010111010100; end
            14'd12884 : begin out <= 64'b1010000011001001101010010110000110101010101011001010010101000100; end
            14'd12885 : begin out <= 64'b1010010011010001001010010100111100101001111101011010001101010000; end
            14'd12886 : begin out <= 64'b0001010001001001101010001100011010100000011011010010010110000101; end
            14'd12887 : begin out <= 64'b1010100010011011001010001100001110101000011000111010101101010011; end
            14'd12888 : begin out <= 64'b1010010001011101101010011101000100101000110111101010000011010001; end
            14'd12889 : begin out <= 64'b1010100101110010001010010100011010101010100001010010011101111010; end
            14'd12890 : begin out <= 64'b0010100011101110101000011110000000101001000100000010100000100100; end
            14'd12891 : begin out <= 64'b1010001001111110100111111100111000100011111011111010101110000001; end
            14'd12892 : begin out <= 64'b0010101100110110101000111000010110101001001010001010010010000001; end
            14'd12893 : begin out <= 64'b0010010011000011101010101101101110101011011101111010100111000100; end
            14'd12894 : begin out <= 64'b0010101010000101101000100101001010101001111001001010001111010001; end
            14'd12895 : begin out <= 64'b0010001000100110101010111001111010101010001011010010101010101111; end
            14'd12896 : begin out <= 64'b0010100001111010101010001111101110101000100010001010101001100101; end
            14'd12897 : begin out <= 64'b0010100010010000101010000100101100011010110110010010101101000101; end
            14'd12898 : begin out <= 64'b0010101100001010001001100010100000101000101010110010011100001101; end
            14'd12899 : begin out <= 64'b0001110110001010101001100110001110101001111111011010100101011011; end
            14'd12900 : begin out <= 64'b1010010100110101101000111001111100100000001110101010101010110010; end
            14'd12901 : begin out <= 64'b0010001010011011001010110111100000101010011010001010100001111011; end
            14'd12902 : begin out <= 64'b1010101100001000100111100001111100100001101111100010011000101000; end
            14'd12903 : begin out <= 64'b1010101010111000101010001100111000101010010001101010101100100010; end
            14'd12904 : begin out <= 64'b0010100001000010000101000011100100101001010001100010100011110101; end
            14'd12905 : begin out <= 64'b1001110110000001001000110000111110100011100011110001111101111001; end
            14'd12906 : begin out <= 64'b0001101011110001101010000110000010100010000111110010101001010010; end
            14'd12907 : begin out <= 64'b0010101111010010001010110010100110101000001000101010100101110110; end
            14'd12908 : begin out <= 64'b1010100011001011001001101011011110101001001110110010001001101011; end
            14'd12909 : begin out <= 64'b1010100010001111101010001000010000101011101010101010010100010010; end
            14'd12910 : begin out <= 64'b1010010100011001101000001111111000100111010010110010100011111100; end
            14'd12911 : begin out <= 64'b1010100000001100001010111100100110101010001101000010011101111101; end
            14'd12912 : begin out <= 64'b1010100101110000001011000100100100100110110011001010001001111010; end
            14'd12913 : begin out <= 64'b1010101111001001101001001101000010101011000100001010100101100010; end
            14'd12914 : begin out <= 64'b1010011100001001001001100000000010101010100011011010101010101011; end
            14'd12915 : begin out <= 64'b0010101000110111101010101001001000100110110011110010100100000001; end
            14'd12916 : begin out <= 64'b1010010000100010101000011110110100100101100010101001100110011001; end
            14'd12917 : begin out <= 64'b1010000111010101001000110111000000101010011010010010100100000110; end
            14'd12918 : begin out <= 64'b0010101100101111001001101011111010100010000011110010010100010110; end
            14'd12919 : begin out <= 64'b1010100101001101001010010101001100100101011000110010101010000101; end
            14'd12920 : begin out <= 64'b1010000101110001001001000001010010100010110001000010100111110000; end
            14'd12921 : begin out <= 64'b1010101011000000101010001001110110101001100101001010100010001001; end
            14'd12922 : begin out <= 64'b1010010101001000001010110010100110100111101000110010001100001001; end
            14'd12923 : begin out <= 64'b1001111000111101101000111011011010100001000000000010100110101001; end
            14'd12924 : begin out <= 64'b1010010010010001101010101001101000100111001101111010101011110100; end
            14'd12925 : begin out <= 64'b1010010001101000100100110001010000101001001000111010001010011101; end
            14'd12926 : begin out <= 64'b0010100110100110101010111111100010100101011101100010000010001100; end
            14'd12927 : begin out <= 64'b0010011011101100001001110100000100100001001000010010100001111011; end
            14'd12928 : begin out <= 64'b0001111100101101001010010001101010101000111000010010101000001110; end
            14'd12929 : begin out <= 64'b1010010101100100001000010010100110100111100101110001111010111101; end
            14'd12930 : begin out <= 64'b0010010000101011000110110000111010010001110000111010110000010100; end
            14'd12931 : begin out <= 64'b1010101011000011001010101001010000100001110111100010010111100110; end
            14'd12932 : begin out <= 64'b1010100111101011001010100111001010101010001111110010011110100101; end
            14'd12933 : begin out <= 64'b1010100100110101001001010110111110001110001101010001101000111111; end
            14'd12934 : begin out <= 64'b0010100100111010000110010100000110100110111001110010001000011011; end
            14'd12935 : begin out <= 64'b1010011000001100101010110110011010100111011010110010101010000110; end
            14'd12936 : begin out <= 64'b0001100110110001001010111010001010101000101010011010001011000001; end
            14'd12937 : begin out <= 64'b1010001101101100001010011110011000101100001100110010001100000001; end
            14'd12938 : begin out <= 64'b1010101101101010001000010100110010011111101110000010100110010110; end
            14'd12939 : begin out <= 64'b1001101111011100101010110101100110100000001000101010000111000001; end
            14'd12940 : begin out <= 64'b1010011101111100101010110001001110101010100000011010101010111101; end
            14'd12941 : begin out <= 64'b1010101010010100001010111101011010101000101000100001100111111100; end
            14'd12942 : begin out <= 64'b0001110101110010001000100010110000100101111101101010011100000000; end
            14'd12943 : begin out <= 64'b1010010110011001101001110100000100101010101001011010101001001101; end
            14'd12944 : begin out <= 64'b0010010011101011101011000000001100101001011010011001111000010000; end
            14'd12945 : begin out <= 64'b1001111000000111101001001001100110011111111010110010011011011111; end
            14'd12946 : begin out <= 64'b0010010100101011101001101101110100101010000111111010010010100111; end
            14'd12947 : begin out <= 64'b0010100110000111001010010010110110101100001111000010101100000101; end
            14'd12948 : begin out <= 64'b0010101011111100101001001110001000101011011001111010100000111111; end
            14'd12949 : begin out <= 64'b0001111111100110101010001101110010100000001111100010100101011111; end
            14'd12950 : begin out <= 64'b1010100111001111101001111010100100100100100000001010011100000100; end
            14'd12951 : begin out <= 64'b1010101100010111100111001011111000101001001000110010101001001011; end
            14'd12952 : begin out <= 64'b1010100010001001101001001101001110011100001111001010101010100010; end
            14'd12953 : begin out <= 64'b0010100010000101101001100001010010011110101101101010101001101110; end
            14'd12954 : begin out <= 64'b0010100111000110001001000101010010100101101001000010101110111101; end
            14'd12955 : begin out <= 64'b0010100100000011100101000110101100100110010101010010011100110011; end
            14'd12956 : begin out <= 64'b0010101110000000001010001011111100100000000111101010100001001010; end
            14'd12957 : begin out <= 64'b0010011110110100101010100111101000101100000100011010100010000101; end
            14'd12958 : begin out <= 64'b1010100011010001101010001011110000101011111001011010010100000001; end
            14'd12959 : begin out <= 64'b1010010110011101001001000010011110100110011101100010011011110010; end
            14'd12960 : begin out <= 64'b1010100101010011001010010010010000101010111111001010101101000111; end
            14'd12961 : begin out <= 64'b0010101010010111101001000010011010010110101001101010011101010010; end
            14'd12962 : begin out <= 64'b0010100110111101101000000000010000100101110000110010010011101010; end
            14'd12963 : begin out <= 64'b0010100101111101101010010110011000011101011101111010010110000100; end
            14'd12964 : begin out <= 64'b1010110000000100101010010010101010101010001001011010011010000011; end
            14'd12965 : begin out <= 64'b1010010010001101001001110110010110100010111011001010100001110000; end
            14'd12966 : begin out <= 64'b0010101011000110001001001110000010010011110100000010101001001001; end
            14'd12967 : begin out <= 64'b1010001010101111001001101000100110100110100100101010011010001001; end
            14'd12968 : begin out <= 64'b0001001011100110001010100100100000100001111101101010010111100010; end
            14'd12969 : begin out <= 64'b1010101111000011001000110000011110101001111110110010101110000110; end
            14'd12970 : begin out <= 64'b0010100100111001100101010001100010100010010101101010100000001101; end
            14'd12971 : begin out <= 64'b1010100011001011001010010000100000100011001011110001110101110000; end
            14'd12972 : begin out <= 64'b1001111011110001001001010001110100101010000000100010011001011111; end
            14'd12973 : begin out <= 64'b0010100111100101001010010000010110100110010011010010000111101101; end
            14'd12974 : begin out <= 64'b1010100001011010100101100011110010100001111011011010010100100000; end
            14'd12975 : begin out <= 64'b0010101101001000001010001000011010101100000010000010101000100001; end
            14'd12976 : begin out <= 64'b1010100101100110101001000101000100101000101111110010010111000100; end
            14'd12977 : begin out <= 64'b0010101001100100101001011000000010100011010010111010100000101011; end
            14'd12978 : begin out <= 64'b1010010011111001101001001100101110100110010111011010100110111111; end
            14'd12979 : begin out <= 64'b0001101011101101001001010000110010011100010100101010100000101001; end
            14'd12980 : begin out <= 64'b1010100100100100101001000000011110011101011101001010100000011111; end
            14'd12981 : begin out <= 64'b0010010011110101101010111101010000100110011001000010101110100101; end
            14'd12982 : begin out <= 64'b0010000110101101101000111011011000011101011011100010101000000001; end
            14'd12983 : begin out <= 64'b0001111101110010101010101111100100011100011001000010100100000011; end
            14'd12984 : begin out <= 64'b1001110000001001001010100000011100100000100110001010101101110010; end
            14'd12985 : begin out <= 64'b1010011110110001001010000011111010101011001110110000000000010101; end
            14'd12986 : begin out <= 64'b0010101001010101001000111100001010101010001111101010000000000101; end
            14'd12987 : begin out <= 64'b1010100000111101001000000111111100101000001000110010100110110101; end
            14'd12988 : begin out <= 64'b1010101110001011001010111101110000101011001011010001000100010100; end
            14'd12989 : begin out <= 64'b1010100000000011101011000000100000101011111000111010011110000001; end
            14'd12990 : begin out <= 64'b0010011101111101001000001000101010100101100000011010101010111101; end
            14'd12991 : begin out <= 64'b1010100001011100001010011110010000100110010010011010101100100111; end
            14'd12992 : begin out <= 64'b0010011001101111101001000111001100101011000000010010011110100000; end
            14'd12993 : begin out <= 64'b1010100110011011101001011111110000101000000111001010011110101011; end
            14'd12994 : begin out <= 64'b0000011011110101101010001101111100100111010100111010001111100110; end
            14'd12995 : begin out <= 64'b1010101001101001101010010101000010101010101111011010010111110000; end
            14'd12996 : begin out <= 64'b1010001011100100000011110110011010101001011001110010100101111000; end
            14'd12997 : begin out <= 64'b0010001111111110101001100110101010100000000101011001110001001011; end
            14'd12998 : begin out <= 64'b1001110011001000101010111110011000100110000100110010100100000111; end
            14'd12999 : begin out <= 64'b0001111110001110001010110100000100101000010010010010010001111010; end
            14'd13000 : begin out <= 64'b1010001001001110101001101111110010101010000010010010101101111010; end
            14'd13001 : begin out <= 64'b1010110000010100000110010110101000101001111101101010010000011111; end
            14'd13002 : begin out <= 64'b0010100000110110001001100111111100100110000000011010100110110010; end
            14'd13003 : begin out <= 64'b1001111011000011100111000100010000101000001000111010011011011100; end
            14'd13004 : begin out <= 64'b0010100011101000101001001010110100101000111000000010100000000011; end
            14'd13005 : begin out <= 64'b0010100000000100101000001100110100100110111011011010101100100111; end
            14'd13006 : begin out <= 64'b0010011001010001101000011111001010100100010001010010100001001011; end
            14'd13007 : begin out <= 64'b0010000101110000001001100011100100100011011011111010100110110110; end
            14'd13008 : begin out <= 64'b0001110010110111100111000000100000101001101001100010101010100111; end
            14'd13009 : begin out <= 64'b0010000111111010101010000100001100100010001111000010101010110100; end
            14'd13010 : begin out <= 64'b0010101011000111001000110010011100101011010100101010011010100010; end
            14'd13011 : begin out <= 64'b1010000100100101101010111001111110101010011001110001111000110010; end
            14'd13012 : begin out <= 64'b1010010101101001101010000101010110101011110101111010011010000001; end
            14'd13013 : begin out <= 64'b1010011010011011001001011110100000101100000110001001011001010001; end
            14'd13014 : begin out <= 64'b0010101011010100100011011011011110101000011110100010101001010010; end
            14'd13015 : begin out <= 64'b0001111101111001101010000101111100100111010110111010100001000001; end
            14'd13016 : begin out <= 64'b1010100010001001000111011111100010101001011010100010101110101111; end
            14'd13017 : begin out <= 64'b0010011101011010001010100111010100100011100011010010010001101001; end
            14'd13018 : begin out <= 64'b1010010101000000001010000011100110101000111010011010101001100101; end
            14'd13019 : begin out <= 64'b1010100100110111101010100000100110100100001000011001110100111000; end
            14'd13020 : begin out <= 64'b0010100110111111101010111001011010100111101011100010010101010011; end
            14'd13021 : begin out <= 64'b0010000101000101101001001001010100101011000100111010000110010001; end
            14'd13022 : begin out <= 64'b1010101100011111101010101001011000101011100000111010000010111111; end
            14'd13023 : begin out <= 64'b1001110011010100001010100110000000101000010110010010001101001011; end
            14'd13024 : begin out <= 64'b0010001110101100001000101011000110101100010100111001101100010000; end
            14'd13025 : begin out <= 64'b0010011011001011001001110010010000100100000010001001101010001110; end
            14'd13026 : begin out <= 64'b1010010111000100000111010110001100100100110010000001110110110110; end
            14'd13027 : begin out <= 64'b0010101000011000001010001001101100011000110000011001101000010101; end
            14'd13028 : begin out <= 64'b0010011100000001100011010011100010001000100011000010010010101000; end
            14'd13029 : begin out <= 64'b1010101000001100001010000101100000100010101000011010100000100101; end
            14'd13030 : begin out <= 64'b1010011010011110001010001001100100101011000001111001101110010101; end
            14'd13031 : begin out <= 64'b1010010110111101101010001000110000011000110100100010100110110101; end
            14'd13032 : begin out <= 64'b1010011110111110101010111001001100101010110101111010101001100001; end
            14'd13033 : begin out <= 64'b0010100001110001101001110110011000100111011001011010011010101101; end
            14'd13034 : begin out <= 64'b0010100111100101001001100010110010011110001001111010101001000001; end
            14'd13035 : begin out <= 64'b1010100001110000101010110101101110101011000000000010011011111011; end
            14'd13036 : begin out <= 64'b1001111000100011101010101011000110101010001000001010100001101111; end
            14'd13037 : begin out <= 64'b1010101101011001001000010101110000100101000100110010000101101010; end
            14'd13038 : begin out <= 64'b1010100001010101101010100111101100100100111010101010100101011000; end
            14'd13039 : begin out <= 64'b0001110110011011001010011101001100100110101001000010011101011100; end
            14'd13040 : begin out <= 64'b1010101000110011001010110000001000101001001100000010100011100011; end
            14'd13041 : begin out <= 64'b0010010110101001101001000111011110011011000000100010101010011100; end
            14'd13042 : begin out <= 64'b1010101110010101001000011010001110101010010101111010100001110110; end
            14'd13043 : begin out <= 64'b0010101100001100001010111001111100011100111001010010000100111000; end
            14'd13044 : begin out <= 64'b1010101101101101001010000110000100100101010011101010101111000000; end
            14'd13045 : begin out <= 64'b0010100111001011001001111100010110100100000111101010101101101011; end
            14'd13046 : begin out <= 64'b1010011100010110001010110010110100101010000100010010101011111100; end
            14'd13047 : begin out <= 64'b1010011010000101101010101000011010101011101000100010100110011011; end
            14'd13048 : begin out <= 64'b1001010011100111001010101011110010101010010110101010011010111101; end
            14'd13049 : begin out <= 64'b1001011001000010001010101101110000100100011011110010100000110010; end
            14'd13050 : begin out <= 64'b1010101100110100001010000010100000100111100111110010010011111000; end
            14'd13051 : begin out <= 64'b0010101011010010000111000101010100100101101100000010101001010001; end
            14'd13052 : begin out <= 64'b0001111010101000101000100110101010100001010011101010100001001101; end
            14'd13053 : begin out <= 64'b0001111010010100101000001001010000011101101100010010011000010100; end
            14'd13054 : begin out <= 64'b0010100100111010001010111011010010100110001000000010100111000111; end
            14'd13055 : begin out <= 64'b0001000011101111001001000000011110101010001111000010011000101000; end
            14'd13056 : begin out <= 64'b1010011001101010101010011110110000100111110101110010100101111100; end
            14'd13057 : begin out <= 64'b1010000010111001001010111101101000101001011010001010001000111010; end
            14'd13058 : begin out <= 64'b0010100000101100001010001001110010100101111011010010011000100010; end
            14'd13059 : begin out <= 64'b0010101100010111001010100001100010100101111000000001101110100000; end
            14'd13060 : begin out <= 64'b0010011100000011101001011111111000100111101110100010011011000010; end
            14'd13061 : begin out <= 64'b1010110000000000000101000011010100100101001011100010100011001101; end
            14'd13062 : begin out <= 64'b0010101100000111101000110010100110101011110001100010101111001011; end
            14'd13063 : begin out <= 64'b0010101110000100001000001010001100101001000010110010100010011110; end
            14'd13064 : begin out <= 64'b0010100000011110101010100011101000100101010111100001110001100110; end
            14'd13065 : begin out <= 64'b0010011011101000101010110100100110101000100101010010010000111101; end
            14'd13066 : begin out <= 64'b1010011000011000000111000010001100101001111000000000101011101101; end
            14'd13067 : begin out <= 64'b1001010011010101101001010110001100100011001111101001101001100011; end
            14'd13068 : begin out <= 64'b1010100000011010001000000101001000100000101010011010010111110110; end
            14'd13069 : begin out <= 64'b0010010110010111101000000011001000101011000111111010011101101100; end
            14'd13070 : begin out <= 64'b0010100010110011101010000000010000101011001011110010101111100100; end
            14'd13071 : begin out <= 64'b0001101101001000101010000000000000100101000101100010100111000110; end
            14'd13072 : begin out <= 64'b1010101100101001101010110011000100100100100111101010100110001110; end
            14'd13073 : begin out <= 64'b0010000010110001101010011010000010100100010010000001000010001110; end
            14'd13074 : begin out <= 64'b0010100101101011000101000011111110100100111010001001000111010000; end
            14'd13075 : begin out <= 64'b0000011111111001101001111100100110100111011110010010100111111000; end
            14'd13076 : begin out <= 64'b0010100010110100101010000000110010101010100000010010100101100000; end
            14'd13077 : begin out <= 64'b1010100100110000100101010001110100100001001111010010010000100111; end
            14'd13078 : begin out <= 64'b0010101110100100000111011000010000100010011111111010101011001111; end
            14'd13079 : begin out <= 64'b0010101101001111101001101101010000100000011110001010100100000100; end
            14'd13080 : begin out <= 64'b1010001011001110101010101101010100011001101110000010100110001111; end
            14'd13081 : begin out <= 64'b0010010100001000100111110110100010100101000110010001011000011000; end
            14'd13082 : begin out <= 64'b0010011000010001101001100001011000101010011100110010100101010010; end
            14'd13083 : begin out <= 64'b0010100010000000101001011110100100100011010101100010101100001000; end
            14'd13084 : begin out <= 64'b1010100011000101100110111011101100010101001111011010000110100001; end
            14'd13085 : begin out <= 64'b1010011010001111000110101111100100101011010000011010010011010110; end
            14'd13086 : begin out <= 64'b0010100010011001001010000110000000101010101011000010011101110001; end
            14'd13087 : begin out <= 64'b1001110110101111000111010010001110011111000101100010000100101111; end
            14'd13088 : begin out <= 64'b1010000101001011001001011010010000100111110101010010010100110000; end
            14'd13089 : begin out <= 64'b0010011101101010101000100111010010101000001011101010101110011000; end
            14'd13090 : begin out <= 64'b1010011101110010001010011011110000100100011101001010101110011011; end
            14'd13091 : begin out <= 64'b0010101011010011101010111011100010100101110111110010100011100011; end
            14'd13092 : begin out <= 64'b1010101011101011101010011100110000101000100001000010101111011010; end
            14'd13093 : begin out <= 64'b0010010011110011001010110011000000101001010111011010101100001101; end
            14'd13094 : begin out <= 64'b1010011111000110101010100101101000101011101010011010101110101111; end
            14'd13095 : begin out <= 64'b0010011101100011101000110001101010100111011010101010100110010111; end
            14'd13096 : begin out <= 64'b1010000110101101001010110110110010100000100100110010000111111101; end
            14'd13097 : begin out <= 64'b0010100100111101001010101100001010101011110011010010101010110100; end
            14'd13098 : begin out <= 64'b1010010101100010101010110000000110100101110001101001101000011001; end
            14'd13099 : begin out <= 64'b0001110001111011101010011000100000101010110111111010001111101111; end
            14'd13100 : begin out <= 64'b0010101100101011101001011100011110101010110001010010010101000011; end
            14'd13101 : begin out <= 64'b1010101100001001001010011100101100100111101111100010001001010010; end
            14'd13102 : begin out <= 64'b0010101000011001101001010010010010101000101110100010100000100010; end
            14'd13103 : begin out <= 64'b1010011100000001001001011110110100100110000001101001100001111111; end
            14'd13104 : begin out <= 64'b1010000111100100001001111001010110101000011001001010011001100101; end
            14'd13105 : begin out <= 64'b0010101100000001001001110111101000101001100001011010000100011101; end
            14'd13106 : begin out <= 64'b0001101110110110100111011000001000101000000000010010101011000111; end
            14'd13107 : begin out <= 64'b1010001000100010101001011000010010100011110001010010101110101101; end
            14'd13108 : begin out <= 64'b0010101001101010001010111011001100010100001011101001100101110010; end
            14'd13109 : begin out <= 64'b1010101001001110100110111100111110101000111011101010010111111110; end
            14'd13110 : begin out <= 64'b0010101011010010001001110101000000101001111100011001100010001111; end
            14'd13111 : begin out <= 64'b1001010000100111001010100111011000101010010010101010000110000000; end
            14'd13112 : begin out <= 64'b0010101100011001001000100001011100101000000101001010010111000110; end
            14'd13113 : begin out <= 64'b1001001111110110001010101011100000010001010111101010010110001011; end
            14'd13114 : begin out <= 64'b1001101110001010101001010010111000101001001111000010010000100101; end
            14'd13115 : begin out <= 64'b0001111010100001001010100010010010100000011010110010011000111110; end
            14'd13116 : begin out <= 64'b0010100100111000101010101010111010101001010000100010010001000101; end
            14'd13117 : begin out <= 64'b0010001000111100100111001110010010100000010100110001011110001111; end
            14'd13118 : begin out <= 64'b1010010100100011001010101000001000100100111100101001110000000010; end
            14'd13119 : begin out <= 64'b0001110111111101101000111011001100100111110011101010010011100010; end
            14'd13120 : begin out <= 64'b0010101111000110101010011000111100101010100110111010010101011100; end
            14'd13121 : begin out <= 64'b0010100000110001101010000001001110100110101110101001110010111001; end
            14'd13122 : begin out <= 64'b1010101110101001001010100111110000101010010001100010100010101110; end
            14'd13123 : begin out <= 64'b1010100111101001100111100000111100100110110101001010101001010111; end
            14'd13124 : begin out <= 64'b0010001100010101101001110111100010101001110001011010010010101101; end
            14'd13125 : begin out <= 64'b0010011111001010101010101100000110101000111111001010101001110000; end
            14'd13126 : begin out <= 64'b0010010100010000000111011100000110101001111111101010100100100010; end
            14'd13127 : begin out <= 64'b0001110100001110100110000111111000100111010001111001011110100000; end
            14'd13128 : begin out <= 64'b0010010101110100001010000011101010100000011000010010100111011001; end
            14'd13129 : begin out <= 64'b0010010110110010001000000101111010101010110100110010001011101110; end
            14'd13130 : begin out <= 64'b1010101011010001101010111101111110101010011010101010100010100001; end
            14'd13131 : begin out <= 64'b1010100101110100001010000110011000011111100001100010010111010110; end
            14'd13132 : begin out <= 64'b1010000100110000001010101100111100101001011001000010011111110001; end
            14'd13133 : begin out <= 64'b0010100110111011001001011011101100101000011101001010000001010000; end
            14'd13134 : begin out <= 64'b0010100110111101001010111010101110100001010110101000110111001100; end
            14'd13135 : begin out <= 64'b1010101000001001101000111111011100101011001010111010010010010111; end
            14'd13136 : begin out <= 64'b1010000111110110001001011111110000101000010011001010000100011000; end
            14'd13137 : begin out <= 64'b0010101010001111101010101011100010100110101011011010101001100110; end
            14'd13138 : begin out <= 64'b1010101100001001001010110001101110101001011100110001111011001100; end
            14'd13139 : begin out <= 64'b1001110111100101101001100011010010100111010100011010100111000011; end
            14'd13140 : begin out <= 64'b0010101101000001101001110111101100101010100001011010011100101001; end
            14'd13141 : begin out <= 64'b0010011011011010000110110111011100101001000111101010010010001101; end
            14'd13142 : begin out <= 64'b0010011100101101001001011011110110100101010101101010101001011011; end
            14'd13143 : begin out <= 64'b0010011100000101001010010111110010101011011001100000100011110110; end
            14'd13144 : begin out <= 64'b0010101001101001001011000000000110101001000010001010010000000010; end
            14'd13145 : begin out <= 64'b1010011001100000001010110000000110101011011000001010101010101110; end
            14'd13146 : begin out <= 64'b0010000101001110101010001011001010100101101001101010001000110000; end
            14'd13147 : begin out <= 64'b0010101100100100001000100000101110101000011001011010101000010011; end
            14'd13148 : begin out <= 64'b1010011001101110101000100101000000101001001101101001111011000001; end
            14'd13149 : begin out <= 64'b0010100010011110101010101011011000100011100110101010000010000101; end
            14'd13150 : begin out <= 64'b1010101110100001101010100011001000101000010001001010000000001001; end
            14'd13151 : begin out <= 64'b1001110100001011101001100101010100101010111011000010100101011001; end
            14'd13152 : begin out <= 64'b0010010110100010101001001011010010101000101101000010010010011011; end
            14'd13153 : begin out <= 64'b1010100000110011000111011100111000101000011100000001101010001101; end
            14'd13154 : begin out <= 64'b1010101001101011000100101011100110100011011001010010100100110011; end
            14'd13155 : begin out <= 64'b1010101000010110001010110101010000101001101001010010101101110110; end
            14'd13156 : begin out <= 64'b0010011101110001101010110011010100100110101011111010101000010100; end
            14'd13157 : begin out <= 64'b1001100101000011101010100111011100011111011001011010011111110100; end
            14'd13158 : begin out <= 64'b0010010011000010101001010011000010100111100101110010011000010100; end
            14'd13159 : begin out <= 64'b0001111011111111001001110110000010101011010010000010011011011111; end
            14'd13160 : begin out <= 64'b0010101001001100001010001010111100101010000101000010101100001111; end
            14'd13161 : begin out <= 64'b0010001111111101101010110100010100100000110001011010101001011101; end
            14'd13162 : begin out <= 64'b1010011110110110001010001000111000101011001011100010100011101001; end
            14'd13163 : begin out <= 64'b0010100111001111101001110000011000011111111011000001110100010110; end
            14'd13164 : begin out <= 64'b1010100000001111101010110101010000011100100001101010001111010101; end
            14'd13165 : begin out <= 64'b0010101000111011101000000111111100101010011000101010001001011011; end
            14'd13166 : begin out <= 64'b1001101010000000101001101111111010100001000110011001110101100000; end
            14'd13167 : begin out <= 64'b1010100100000010101010100000110110011010110010011010011001010010; end
            14'd13168 : begin out <= 64'b1010101101111000101010111101011110101000110110111001110010001010; end
            14'd13169 : begin out <= 64'b1010011101100010101010100000111010101001111001110010100101010001; end
            14'd13170 : begin out <= 64'b0010100100001100001001100101010000100011011010111010101011000011; end
            14'd13171 : begin out <= 64'b0010101011101111101000000000110100100101111100101010000100101101; end
            14'd13172 : begin out <= 64'b0010100100100110001010111011111000100110100100000010100110110101; end
            14'd13173 : begin out <= 64'b1010100011000011001010010111101000101011001000010010011001001000; end
            14'd13174 : begin out <= 64'b0001011101101101000111111111010010100000111000101010010100111100; end
            14'd13175 : begin out <= 64'b1010000000110111001010010111100000100100001100101010101001000001; end
            14'd13176 : begin out <= 64'b1010001000110001101010011100100010011110001000001010101111001001; end
            14'd13177 : begin out <= 64'b1010011101011110101001111011001110101000000100101010100110011010; end
            14'd13178 : begin out <= 64'b1010010001100001101001110000101010100110111010011010010111100100; end
            14'd13179 : begin out <= 64'b0001100100000000001010011110101010100100110101100010101100100011; end
            14'd13180 : begin out <= 64'b1001100101010111001010000110110010101000001010100001110000000011; end
            14'd13181 : begin out <= 64'b1010010011110000001010010011000100100100111100110010100000010111; end
            14'd13182 : begin out <= 64'b0001110001100100101001010110011000101001111110001010100111000011; end
            14'd13183 : begin out <= 64'b1010101011111000101010001001100110101010010111010010100000000111; end
            14'd13184 : begin out <= 64'b1010011101100001101010010111001000100100111011110010100101110100; end
            14'd13185 : begin out <= 64'b1010011010000110101000001010100010101010100100000010100100100010; end
            14'd13186 : begin out <= 64'b0010000100101101101001110011010000101001101000100010100001000000; end
            14'd13187 : begin out <= 64'b0000000111010001100101010110001000100101100001000010100100010111; end
            14'd13188 : begin out <= 64'b0010101101100011001010110000100010100000110110110010101111011011; end
            14'd13189 : begin out <= 64'b1010100111101011101010110101101100100101011110010010101010111101; end
            14'd13190 : begin out <= 64'b0010100110101001100101111011110110101011011110110010100011111000; end
            14'd13191 : begin out <= 64'b0010000011101010101001000000001100100101010010001001110110011110; end
            14'd13192 : begin out <= 64'b1010100011101011001010001110110010100011001100110010100111010000; end
            14'd13193 : begin out <= 64'b1010101000001010101010100011001010101011011011000010100111000100; end
            14'd13194 : begin out <= 64'b1010100001011110001001000111000100101011011010010010100100101100; end
            14'd13195 : begin out <= 64'b1010101011011000001010011111111110101001000100100010100111010000; end
            14'd13196 : begin out <= 64'b0010010000110011101001101100111110100001011011100010101111000101; end
            14'd13197 : begin out <= 64'b1010001000011000001010011101101110100111010101010010001110100111; end
            14'd13198 : begin out <= 64'b1010100011101101101010111111110100100010100000111010100000110111; end
            14'd13199 : begin out <= 64'b0010101110001110001010010101011010100100101100110010010000010101; end
            14'd13200 : begin out <= 64'b1010101011110100101010101100101110101011101011011000110001010001; end
            14'd13201 : begin out <= 64'b0010101001001000101010000101000000101001100110010010011010100111; end
            14'd13202 : begin out <= 64'b1010011110010011001001000110101100101001111110110010011101001110; end
            14'd13203 : begin out <= 64'b0010101100101001101010000001001010100100001011010010001111011110; end
            14'd13204 : begin out <= 64'b0010100100111111001010101000001100011000001101000010000100010110; end
            14'd13205 : begin out <= 64'b1010011000111100001010011110110100100101001001111010100000100111; end
            14'd13206 : begin out <= 64'b0001100011001110000111101110101110101011011100110010100001110101; end
            14'd13207 : begin out <= 64'b0010100001100100101001001101110000101001000100011010100011011111; end
            14'd13208 : begin out <= 64'b1001110101001111001010010100100100100011110011010010101001010111; end
            14'd13209 : begin out <= 64'b1010010101100001000100001000001000101011110000100010010011001101; end
            14'd13210 : begin out <= 64'b1010001011100011000110111110111100101001011101101010011001010101; end
            14'd13211 : begin out <= 64'b1001011010000101101001001100101010101010110111011010101000100110; end
            14'd13212 : begin out <= 64'b1010010000010000001001011110101110101000110010101010011101100010; end
            14'd13213 : begin out <= 64'b1010000100011101001010111001001100101010001011000010101100100000; end
            14'd13214 : begin out <= 64'b0010001111010000000111101110111100100011100100000010001010010111; end
            14'd13215 : begin out <= 64'b0010100001000011101001010100111110101001001001101001110010101100; end
            14'd13216 : begin out <= 64'b0010101001100110001010110011101110101001010010101010001000011101; end
            14'd13217 : begin out <= 64'b0010100111101110101010111001110000100100101101000010011101000100; end
            14'd13218 : begin out <= 64'b0010100111000111001001101101101110100111101001011010100000001000; end
            14'd13219 : begin out <= 64'b0010100100001000001010100011000100100011111101111010000111110111; end
            14'd13220 : begin out <= 64'b0010101110001001101001110000001010011001100011111010011110001100; end
            14'd13221 : begin out <= 64'b1010100111001100001010111010101010101001000011101010001001011111; end
            14'd13222 : begin out <= 64'b0010100110010110001000100100011110101000000010110010100111110010; end
            14'd13223 : begin out <= 64'b1010010001011001001010111110000010011000101111100001101001100101; end
            14'd13224 : begin out <= 64'b1010101000111101101001110011111010100100010010000010101010010100; end
            14'd13225 : begin out <= 64'b0010010100010001101001110111110010101010111101101010000110011001; end
            14'd13226 : begin out <= 64'b0010101000001101001010011010011000100010110011011010100011010010; end
            14'd13227 : begin out <= 64'b0001111001000001101010110100101010100100010100010001111101001111; end
            14'd13228 : begin out <= 64'b1010100001111001001001001100110010101000000010001010101011101010; end
            14'd13229 : begin out <= 64'b0001110000111100001001001100000110100001011000000010100101000010; end
            14'd13230 : begin out <= 64'b1010100001000100101010011110110110101000011111110010011000011010; end
            14'd13231 : begin out <= 64'b0010100000011110101010011010010010101000010110010001001111100010; end
            14'd13232 : begin out <= 64'b0010100001000111101001010000101100101011101110100010010000100101; end
            14'd13233 : begin out <= 64'b1010100011010000101010010101110110101000010010111010011001001001; end
            14'd13234 : begin out <= 64'b1010101011100000101010110111001000101000111110110010011111000111; end
            14'd13235 : begin out <= 64'b0010101101110100100111010100001000101000010100011010010100110110; end
            14'd13236 : begin out <= 64'b1010101101101011001001000001010010100000011010110010011001010010; end
            14'd13237 : begin out <= 64'b0010101011111010101000001111000110101001100100100010001100111111; end
            14'd13238 : begin out <= 64'b1010101010011000000111110100000110100111110100010001100100011001; end
            14'd13239 : begin out <= 64'b0010101101101100101010000001001100101001111110001001011001111001; end
            14'd13240 : begin out <= 64'b0010101011010010101010011100011010011011100110000010010110110010; end
            14'd13241 : begin out <= 64'b0010101110111000001010110111101100100100001101000010101001000001; end
            14'd13242 : begin out <= 64'b1010011011111100101010001001000100101010001101010010011100000100; end
            14'd13243 : begin out <= 64'b0010101100101000001001001111011000101010000100110010101011011000; end
            14'd13244 : begin out <= 64'b0010100110000111101010011001111000100110000011100010101110101011; end
            14'd13245 : begin out <= 64'b1010010100011011001000000011100010101011000011010001001111010110; end
            14'd13246 : begin out <= 64'b0010010110001111101010101000011010100011011101110010101111010100; end
            14'd13247 : begin out <= 64'b1010101011001111101000100110110010101010001110001010100010010010; end
            14'd13248 : begin out <= 64'b1001110010101001100111101100001100100000000110111000111111000010; end
            14'd13249 : begin out <= 64'b0001010111110000101000010101010110100101011010111010101110011111; end
            14'd13250 : begin out <= 64'b1010101110000101001010100111110100100000001110000010101000101111; end
            14'd13251 : begin out <= 64'b1000110110010000001010100000110100010000100101010010101111000000; end
            14'd13252 : begin out <= 64'b0010010110010100000101111111011010100100001001001010101110001010; end
            14'd13253 : begin out <= 64'b1001110001001010001010000011110100100000110011101010001110000000; end
            14'd13254 : begin out <= 64'b1010100000111010001001001010011100100110110000001010101000110110; end
            14'd13255 : begin out <= 64'b1010100101001010000110111101011000100011111110010010011011101110; end
            14'd13256 : begin out <= 64'b0001101011010110000001010011010010101010101101000001111101100000; end
            14'd13257 : begin out <= 64'b1010001001110001100111110100001110100011011101101010010100011111; end
            14'd13258 : begin out <= 64'b1010101011111000000111000000100110010011110110011010100110011001; end
            14'd13259 : begin out <= 64'b0010001001011011000100100010010100101010110111101010101001010010; end
            14'd13260 : begin out <= 64'b1010101101100000001001010101011010100101011101101010100111001000; end
            14'd13261 : begin out <= 64'b1001100011101011001010010011101100100110100101101010011011011110; end
            14'd13262 : begin out <= 64'b0010100100110100001001011000001010100111101011001010010010111111; end
            14'd13263 : begin out <= 64'b1010011010100001001010011010001110100110100100101010101111001101; end
            14'd13264 : begin out <= 64'b0010101111100010101001101001101110101001101000110010100111111000; end
            14'd13265 : begin out <= 64'b0010100010101100001010100001011010101001010011110010010111010101; end
            14'd13266 : begin out <= 64'b0010001100011111101010000011111110100111111110001010101001100010; end
            14'd13267 : begin out <= 64'b1010100101101101101000011100000100100010100111001010000110101000; end
            14'd13268 : begin out <= 64'b0010101000011000001010100100100100101011000000001010101100101001; end
            14'd13269 : begin out <= 64'b0010010000100111001001111000101000101010111001011010011111010110; end
            14'd13270 : begin out <= 64'b0010101100111100101010010000110000010111111111001010100111011000; end
            14'd13271 : begin out <= 64'b1010101011010100101000011101110110011011110101001010100001001001; end
            14'd13272 : begin out <= 64'b0001100111001110001010001100000100100110000101000010010101110001; end
            14'd13273 : begin out <= 64'b0010100011010111001000010100111010101010000000110010010010111011; end
            14'd13274 : begin out <= 64'b1010101100100000101001010101111100100001100001100010011011001001; end
            14'd13275 : begin out <= 64'b0010010000011001101000100000010100100100000011110010101101010000; end
            14'd13276 : begin out <= 64'b0001110110101100001001011101001010011100100101110010001111110010; end
            14'd13277 : begin out <= 64'b0010010000101001001010000100000100100100001111100010010001000011; end
            14'd13278 : begin out <= 64'b0010100101110111101010110111011010100110100001010010100001010010; end
            14'd13279 : begin out <= 64'b0010100001101101101001110101000000100111001101100001001100000010; end
            14'd13280 : begin out <= 64'b0010011000110001001001000111101110101011011010001010101110110000; end
            14'd13281 : begin out <= 64'b0010110000111000001000001011000010100111100110101010101101111110; end
            14'd13282 : begin out <= 64'b1010010000011110101010101110010100101000011101111010101011100000; end
            14'd13283 : begin out <= 64'b1010000011010010001010100101011000100001111000010010100011010110; end
            14'd13284 : begin out <= 64'b0010100000100010101001111101001000100110010011111010011011010001; end
            14'd13285 : begin out <= 64'b1010100011011111101010110001001000101010000001100010101111001101; end
            14'd13286 : begin out <= 64'b1010100001010101001010111001011010100010110110001010001101001000; end
            14'd13287 : begin out <= 64'b1010101101011010101000001011001000101010111011100001011101011011; end
            14'd13288 : begin out <= 64'b1010101110100101001000000011011100100011111110110010010101110001; end
            14'd13289 : begin out <= 64'b1010100100101101101001101011011110101010110110110010101101110111; end
            14'd13290 : begin out <= 64'b0010011110011010001001110011100010100101101110001001010011101111; end
            14'd13291 : begin out <= 64'b1010100110001000001010110001101100101011101011100001001011101001; end
            14'd13292 : begin out <= 64'b0010101100100000001001011100001100101000100001010010101011110111; end
            14'd13293 : begin out <= 64'b1010101111010010001010110100110100100000110111010010100000111101; end
            14'd13294 : begin out <= 64'b0010011001101010001000000110011110011100010001111010001011010001; end
            14'd13295 : begin out <= 64'b1010001010110000001010011010100000100011111001100000010011010110; end
            14'd13296 : begin out <= 64'b1010101101001000001000111101001100101001010000010010101111100110; end
            14'd13297 : begin out <= 64'b0010000100010100001000101110010100101000100011110010100100101111; end
            14'd13298 : begin out <= 64'b1010001111000100101010011011010110100110011110000010100101010111; end
            14'd13299 : begin out <= 64'b1010001100010000101010110010100000100101110001101010000010011001; end
            14'd13300 : begin out <= 64'b0010011111011010000111001010001010101010110000001001001011111010; end
            14'd13301 : begin out <= 64'b0010100011000001000110011011110100100110011110101001111111100110; end
            14'd13302 : begin out <= 64'b0010100110101111101010100110011110011010001000001010100110111101; end
            14'd13303 : begin out <= 64'b1001011000000110001001010100010010101010111001110010010001011110; end
            14'd13304 : begin out <= 64'b1010001000100111001010010111010110101000100011001010001111001101; end
            14'd13305 : begin out <= 64'b1010100111001111001001111011101000100111001010111010101001100000; end
            14'd13306 : begin out <= 64'b0010101100001000101010001000100010010001101011100010001100100110; end
            14'd13307 : begin out <= 64'b0010101100101001001001010101100010100001000101001010001101111001; end
            14'd13308 : begin out <= 64'b0010011010111001001010100010101100100101010000101010101111110100; end
            14'd13309 : begin out <= 64'b0010100001110000001010001100011100101000000010010010100011111110; end
            14'd13310 : begin out <= 64'b1010101001000111101010110100110010100011100011100010101010100101; end
            14'd13311 : begin out <= 64'b1010101100000000101010011010010100101001001100011010000000011111; end
            14'd13312 : begin out <= 64'b1010001000001011001000010001110110100111000111100010101001011011; end
            14'd13313 : begin out <= 64'b1010100001010100001001110011000100101011100011111010100111011000; end
            14'd13314 : begin out <= 64'b1010101000000000101010010000101000101000010000100001001011110100; end
            14'd13315 : begin out <= 64'b1010101100101111000110110110100000100010110101011010010100101100; end
            14'd13316 : begin out <= 64'b0010100001011000101000101011100110101001100001011001100011110100; end
            14'd13317 : begin out <= 64'b1010010111111010000111111010101000101011001000001010001100010100; end
            14'd13318 : begin out <= 64'b1010101011000001101010010100100110101001101111100010001111101110; end
            14'd13319 : begin out <= 64'b0010100000010011101010010000001100100000101001100010010111101111; end
            14'd13320 : begin out <= 64'b0010011101111010101000111001100000101011011011000010011111010111; end
            14'd13321 : begin out <= 64'b0001111000001011000110001000110110100101110101110010000010000111; end
            14'd13322 : begin out <= 64'b1010010101110101101001011000111000101001100001100010010001001101; end
            14'd13323 : begin out <= 64'b1010100001001001001010101001011000101000011010000010100010101101; end
            14'd13324 : begin out <= 64'b1010101100101101001010101001000010101001010110110001101111110111; end
            14'd13325 : begin out <= 64'b1010001011100010101010101000110010101011111110111010001100010100; end
            14'd13326 : begin out <= 64'b1010101011101011001010001110111010100111110000110010011111000100; end
            14'd13327 : begin out <= 64'b0010001101100111001010100100010010101000001001110010101001001000; end
            14'd13328 : begin out <= 64'b1010011000101110001010111110010010101010011111100010101011000000; end
            14'd13329 : begin out <= 64'b1010011111010001100110100001100010010010111111001010101111011111; end
            14'd13330 : begin out <= 64'b1010011111110101101001000110001110100100111110100010101010111111; end
            14'd13331 : begin out <= 64'b1010100010111100101010110101011000101011111110100010011111000100; end
            14'd13332 : begin out <= 64'b1010101100000000100111100110000110100101110110111010011111100110; end
            14'd13333 : begin out <= 64'b0010101101000000001001010110011010101010111000100010100110101100; end
            14'd13334 : begin out <= 64'b0010100100001110001000111110110100100111011011100010101010000001; end
            14'd13335 : begin out <= 64'b0010011010010011001001111001101010101011101111000000100101010011; end
            14'd13336 : begin out <= 64'b1010101101001011001000011100011100011110011110000010010000101010; end
            14'd13337 : begin out <= 64'b0010100000010111001010010111000010100100111001001010100010000100; end
            14'd13338 : begin out <= 64'b1001101111000010101001110001001100101010101110001010100100001011; end
            14'd13339 : begin out <= 64'b1010001010001110001001001001010100001110101101100010011000010001; end
            14'd13340 : begin out <= 64'b0010100001100000101001101010100000101011111100011010011001011100; end
            14'd13341 : begin out <= 64'b0010001111011101001010110000011000101010010111110010101001101111; end
            14'd13342 : begin out <= 64'b0010010001000101001001011001010000101000111110110010000001010000; end
            14'd13343 : begin out <= 64'b0010101000001000001010000111000110101010010101100010010110010010; end
            14'd13344 : begin out <= 64'b0010100101100011101010001010011000101010110001101001111100110100; end
            14'd13345 : begin out <= 64'b0010011010100011100101100000110100100101000001010010010001100010; end
            14'd13346 : begin out <= 64'b0010100000100000001001001100100100011010110001100010010100011111; end
            14'd13347 : begin out <= 64'b0000110000101010101000100101011000100001011100011010100100111000; end
            14'd13348 : begin out <= 64'b1010011001101001101010100001111000101011100010100010101010011001; end
            14'd13349 : begin out <= 64'b0001100000111100001000100101110110100100110001110010101001010100; end
            14'd13350 : begin out <= 64'b0010100010101010101001110111001010100101010101000010100000100011; end
            14'd13351 : begin out <= 64'b0001110011001011101001001010111000011000101111111010011101000101; end
            14'd13352 : begin out <= 64'b1010101100110111001001010000011100100011010100100010100000110001; end
            14'd13353 : begin out <= 64'b0010011100001010001010100101100000101010011111111010001110000000; end
            14'd13354 : begin out <= 64'b1001100011000011101001101101111100100111011001100010101011111010; end
            14'd13355 : begin out <= 64'b1010001000011111101001011011110100100101110000011010011001000101; end
            14'd13356 : begin out <= 64'b0010100001100100001010011001110100101001001100111010101000001011; end
            14'd13357 : begin out <= 64'b0010011101010001001010001101110000100100110001010010101011111011; end
            14'd13358 : begin out <= 64'b1010100110010100001010011111100000100111111111000001111001010111; end
            14'd13359 : begin out <= 64'b0010100010011110101010101111010110011101010101111010011000101111; end
            14'd13360 : begin out <= 64'b0010011100001011001001010010100000101000010011011010101111111011; end
            14'd13361 : begin out <= 64'b0010101111100100101010110111100010101000000011010010101110111111; end
            14'd13362 : begin out <= 64'b1010010110001100101001011011010100101001100111010010101001111101; end
            14'd13363 : begin out <= 64'b1010100001011100001010111101101010100111110111011010101010101011; end
            14'd13364 : begin out <= 64'b0010001001011010100111111000100110101001101001101010100001011001; end
            14'd13365 : begin out <= 64'b0010101111001011000111110111000100100011101010100010000101011101; end
            14'd13366 : begin out <= 64'b0010100001001010001000000110011110101011010110101010101000010011; end
            14'd13367 : begin out <= 64'b0010010010000110001001111100010000101010101001110010100101110111; end
            14'd13368 : begin out <= 64'b1010010010101010001010000101010000011011000111001010011001100100; end
            14'd13369 : begin out <= 64'b0010001101010001001001100100010110101000100100110001011101111000; end
            14'd13370 : begin out <= 64'b1010100110100100101010101100100000100010111111010001101111100001; end
            14'd13371 : begin out <= 64'b1010100011010010101001110110101110101010111010011001101101101000; end
            14'd13372 : begin out <= 64'b0010100010100011001000011101000010011100001101110010101100111000; end
            14'd13373 : begin out <= 64'b0010011010101111001010110110001000011100100110001010101011011110; end
            14'd13374 : begin out <= 64'b0010000011100110101010000000110110100001010001010010010011011001; end
            14'd13375 : begin out <= 64'b0010010001000010101010001010010110101001000011001010101110001000; end
            14'd13376 : begin out <= 64'b1010010010100000100110011100010100011000011011100010101010111001; end
            14'd13377 : begin out <= 64'b0001111000011011101010010101101000101011010111000010100000100001; end
            14'd13378 : begin out <= 64'b1010100000011010001010000011110100100111001000101001111101011110; end
            14'd13379 : begin out <= 64'b0010011110000111000111010000010000011001100110001010001010100000; end
            14'd13380 : begin out <= 64'b1010101001100110101001101100000000101011101000000001110011000010; end
            14'd13381 : begin out <= 64'b1010011001111010101001101010000110101010110010010010011111101101; end
            14'd13382 : begin out <= 64'b1010010101000101001001101011111000101011011110101010010001011001; end
            14'd13383 : begin out <= 64'b0001000010110000001000010100011010011110100101110001101100110010; end
            14'd13384 : begin out <= 64'b1010010110011110001010100111011110101011000011111010100110111100; end
            14'd13385 : begin out <= 64'b1001011100001011100110011100100100101011101001010010011011110010; end
            14'd13386 : begin out <= 64'b1010101100011011001000011100000100101010111010101010101011011010; end
            14'd13387 : begin out <= 64'b1010101110000111001010010010000010101010111101100010100101110011; end
            14'd13388 : begin out <= 64'b1010101011111011001010011011110100101001011001100010100111110001; end
            14'd13389 : begin out <= 64'b0010100000101111001001110000110000100001101011111010001010001010; end
            14'd13390 : begin out <= 64'b1010110000000001101010101100000110101010100100111010101011100010; end
            14'd13391 : begin out <= 64'b1010100001011111101001011101011100100101100000101001111010100100; end
            14'd13392 : begin out <= 64'b0010100100001100101001011001100100101000011100001001010001000010; end
            14'd13393 : begin out <= 64'b0010100010101100101010101111100110100101100111111010100110001111; end
            14'd13394 : begin out <= 64'b1010100000110111101000011001111010101001011010111010101110000100; end
            14'd13395 : begin out <= 64'b0010011111111111101001100000111110100111111100001010011000110011; end
            14'd13396 : begin out <= 64'b1010011011110101100111110110010100100101101011110010011000000100; end
            14'd13397 : begin out <= 64'b1010001010110001001010100110110000100100101011010010000000000001; end
            14'd13398 : begin out <= 64'b0010000000001100101001100011101000100111001011000010101001100000; end
            14'd13399 : begin out <= 64'b0010011010011011101010010001011000100011010010111001111000011001; end
            14'd13400 : begin out <= 64'b1010100011111100000111111110111000101011011111010010100111001000; end
            14'd13401 : begin out <= 64'b1010101101101100101010010001010100100101011001010001001011111010; end
            14'd13402 : begin out <= 64'b1010101001010100100110100100110000101010000100000010101010000001; end
            14'd13403 : begin out <= 64'b0010100100100101101000011101010010100101000111110010101000001111; end
            14'd13404 : begin out <= 64'b0010100101101011000110010001010100011011000010001010001111110111; end
            14'd13405 : begin out <= 64'b0001100001010110101000010001110110100110011000100010101111101001; end
            14'd13406 : begin out <= 64'b1010011001010001101010001000010110100111110000101010100001111000; end
            14'd13407 : begin out <= 64'b0010011011101000001010010100111010101011110010001010011001100111; end
            14'd13408 : begin out <= 64'b1010100010100010101000000110011010101001101000101010100100011100; end
            14'd13409 : begin out <= 64'b0010100010011000101001001100000010100101100110110010101000101100; end
            14'd13410 : begin out <= 64'b0010011100000100101010001011000010101010000111100010100110011011; end
            14'd13411 : begin out <= 64'b0010101001000110101001011001100110101001110000000010100000001111; end
            14'd13412 : begin out <= 64'b0010101110110001001001011010101010101011110111010010101011010111; end
            14'd13413 : begin out <= 64'b1001110011011100001000011100011010100000011011110010100001110111; end
            14'd13414 : begin out <= 64'b0010000100000000101010000010101000100010000101101010010001111011; end
            14'd13415 : begin out <= 64'b0010010101111011001000000111110000100101010011110010100101110111; end
            14'd13416 : begin out <= 64'b0010001101101111101001110001010010011111101011101010100000110111; end
            14'd13417 : begin out <= 64'b1010101110010001101010001011111100011101000110010001111100101000; end
            14'd13418 : begin out <= 64'b1010100111010110001010111011011110100001110001000010000101000000; end
            14'd13419 : begin out <= 64'b0010100101111000001010110001111010101011101101000010101100101100; end
            14'd13420 : begin out <= 64'b1010101001101000101010001101011000100010101100001001111011000010; end
            14'd13421 : begin out <= 64'b1010100001101110001001001010101110101001110010111010010110001011; end
            14'd13422 : begin out <= 64'b1010010100101101001010101001011110011011000001110010101101101000; end
            14'd13423 : begin out <= 64'b0010100110011110101010001000101010011110001100110010101011000010; end
            14'd13424 : begin out <= 64'b0010011101001010101010111001110100101000100011101010101111100011; end
            14'd13425 : begin out <= 64'b1010100100010111101010010011100000100110000011111010011101110011; end
            14'd13426 : begin out <= 64'b1010100101011111001010000000001100100001000101110010100000111000; end
            14'd13427 : begin out <= 64'b0001010001011111101001001001001010101000111011100010101001100111; end
            14'd13428 : begin out <= 64'b1001101011111001001010111010111100101001011110001010011111111011; end
            14'd13429 : begin out <= 64'b1010000111100100001000001010100100101001001100011010010111101110; end
            14'd13430 : begin out <= 64'b1010001000000000100101110001100010100111010110010010100011100111; end
            14'd13431 : begin out <= 64'b0010000001101100001000100001110100010100100000011001011001111111; end
            14'd13432 : begin out <= 64'b0010010011011110001001010011011000100011001000110010101101101010; end
            14'd13433 : begin out <= 64'b1010100010101010000111100011001010011101100011101010101101110001; end
            14'd13434 : begin out <= 64'b1010101000001011001010101100110100011000010011011010100100111001; end
            14'd13435 : begin out <= 64'b1001011011110100100111010101111010101001110011111010100001001011; end
            14'd13436 : begin out <= 64'b0010100010010100101001100001000000100011101000101010101001010111; end
            14'd13437 : begin out <= 64'b1001111111100011101010001000101110100111101110110010101110110000; end
            14'd13438 : begin out <= 64'b0010000010011011101010010000101000011001110001010010011101111000; end
            14'd13439 : begin out <= 64'b0010101100111101100101110100110010011010100111100010101101111010; end
            14'd13440 : begin out <= 64'b1010011011101010101010100010001100101011010010001010010001101011; end
            14'd13441 : begin out <= 64'b0010101011010011100111110000011010101011000001001001010110000110; end
            14'd13442 : begin out <= 64'b1010101101100001101010110010011000100100101010011010101100011100; end
            14'd13443 : begin out <= 64'b0010001110001101001001100110100100101000011000100010010001110001; end
            14'd13444 : begin out <= 64'b0010101001110001101001100101011100100100100111101010101010111101; end
            14'd13445 : begin out <= 64'b0010001011001001100011101001110100101011100000010010010111110101; end
            14'd13446 : begin out <= 64'b1010101100100101101010110000111100011101110111101001101000000110; end
            14'd13447 : begin out <= 64'b0001110100110101001010100010111110101010001101000010010111110101; end
            14'd13448 : begin out <= 64'b1010011010111010101001011000100110100100010001111010010100110101; end
            14'd13449 : begin out <= 64'b1010011001010111001010001000001100101011001011101010101101011000; end
            14'd13450 : begin out <= 64'b0010100010101100101001110101111010101010110010000010100000110011; end
            14'd13451 : begin out <= 64'b1001111101110001001010111010110010100001101000110010010100101001; end
            14'd13452 : begin out <= 64'b1010100001011100001010100011000010100000011011100010011001000001; end
            14'd13453 : begin out <= 64'b0010000110010011101001101011010000101010001111110010100010000011; end
            14'd13454 : begin out <= 64'b1001110101100110001001101101000110100001111010101001100011111110; end
            14'd13455 : begin out <= 64'b1010010100111001101001000001010000101010010011001010010110011110; end
            14'd13456 : begin out <= 64'b0010010011110001101010010010000100100111011100001010011110110101; end
            14'd13457 : begin out <= 64'b0010101001111001101001001101010100100011100000101010011111100001; end
            14'd13458 : begin out <= 64'b0010100001011011101010000011011010100101000100011010101101101100; end
            14'd13459 : begin out <= 64'b1010000100000110101010101101110000011100001001000010011010000110; end
            14'd13460 : begin out <= 64'b1010100011111101001010111011101010011000011010000010100100011010; end
            14'd13461 : begin out <= 64'b0010100101011000101000110011101100101001001100111010010110001001; end
            14'd13462 : begin out <= 64'b0010011010000110001001001110010110101011001110111010100011111001; end
            14'd13463 : begin out <= 64'b0010100000011010101010110110110100101000001110000010010011010010; end
            14'd13464 : begin out <= 64'b0010010100101011101001100111110100101010100011110010100001101011; end
            14'd13465 : begin out <= 64'b0001111011000111101010001000101000101001111110010010100111100011; end
            14'd13466 : begin out <= 64'b0001111111000010101010011110010100101000010001011010100101110000; end
            14'd13467 : begin out <= 64'b1010100011110010101000111101001100101011000100110010100100010100; end
            14'd13468 : begin out <= 64'b1010011001100101001010011110011100011110110000100010101000001100; end
            14'd13469 : begin out <= 64'b1010100110101100100111100111010010101011110111010010001001111000; end
            14'd13470 : begin out <= 64'b1010100100110000001001100110000010101000000000001010101101011010; end
            14'd13471 : begin out <= 64'b1010100000011001101010101010101110100100011100010010101100010111; end
            14'd13472 : begin out <= 64'b1010100011010010001010110000101100100100101001001010010101010101; end
            14'd13473 : begin out <= 64'b0010100101001011001001001000111100101000111110011010100011111001; end
            14'd13474 : begin out <= 64'b0010001001010001001010010010111000011110001000001010100001101111; end
            14'd13475 : begin out <= 64'b0010000010011001101010011100111100100110011001001010101111000111; end
            14'd13476 : begin out <= 64'b1010101011110010001010101110010010010100100000000010010100011000; end
            14'd13477 : begin out <= 64'b1010001001000100101010000110001110101010110011010010000011011000; end
            14'd13478 : begin out <= 64'b1010011100101101001001011111111000100100111101100010011011011101; end
            14'd13479 : begin out <= 64'b1010001100010101001010101101011010011101001100101010100000100110; end
            14'd13480 : begin out <= 64'b0010011010000011100110111111101100101000100110001010010011100000; end
            14'd13481 : begin out <= 64'b0010010100010110001010101011101100101001100001100010101010110010; end
            14'd13482 : begin out <= 64'b0010001111111101101001001001100110101011010111010010001100000010; end
            14'd13483 : begin out <= 64'b1001110101001010100110110000110110100100111100101010100000111110; end
            14'd13484 : begin out <= 64'b1010011011001100001010001001010110101011011010011010100011011101; end
            14'd13485 : begin out <= 64'b1010101100101100100111000100111000101011111110000010011010101001; end
            14'd13486 : begin out <= 64'b1010100010111110101010010000000000101010001100000010101111001110; end
            14'd13487 : begin out <= 64'b1001110110001101001010101110110100011111001011111001010010010011; end
            14'd13488 : begin out <= 64'b1010011011110111101000011101011000011111011110110010000010010111; end
            14'd13489 : begin out <= 64'b0010101100110000001010100010110000101011111110000010100101100000; end
            14'd13490 : begin out <= 64'b1010100000011001101001011100001110101001100011100010101110011101; end
            14'd13491 : begin out <= 64'b1010100010101001001000011001110110100001011111111010101110010001; end
            14'd13492 : begin out <= 64'b1010101101001111101000011011011100100011010000100010101100001101; end
            14'd13493 : begin out <= 64'b1010101000011100001010011011111100101001001111011010011000001010; end
            14'd13494 : begin out <= 64'b0010011100111011101000101010000110100010100101000010010100100000; end
            14'd13495 : begin out <= 64'b1010100110100111101010101001010110101010011110000001110100011011; end
            14'd13496 : begin out <= 64'b0010101111101000101010101010000010100111011110100010100001100001; end
            14'd13497 : begin out <= 64'b0001100110001011001001001011110110100101100111111010101001111111; end
            14'd13498 : begin out <= 64'b1010010111110001101000111010101110101000110010100010001001101001; end
            14'd13499 : begin out <= 64'b1010101110000000001000011011101000100111111100101001100000010101; end
            14'd13500 : begin out <= 64'b0010010101000111001001011011100010100011010101010010011110010100; end
            14'd13501 : begin out <= 64'b0010010101001111001000010011011010101001100100011001001100000001; end
            14'd13502 : begin out <= 64'b0010001101010011101010010011001100101000100100110010101000101100; end
            14'd13503 : begin out <= 64'b1010101011000010001001111010010110101000010010011010010101101011; end
            14'd13504 : begin out <= 64'b1010011100110110001001011110101000011101111000101001111101110101; end
            14'd13505 : begin out <= 64'b1010101100100110001000011100011000101011000111001010101100011001; end
            14'd13506 : begin out <= 64'b0010011001011101001001010100010100101001100111101001011111011000; end
            14'd13507 : begin out <= 64'b1010001001100100001000110100110000011111100101101010001011010111; end
            14'd13508 : begin out <= 64'b0010101010100001100001100001010000101001111111111010001101111110; end
            14'd13509 : begin out <= 64'b1010101000001001100100011000110110011101100010111010000010101100; end
            14'd13510 : begin out <= 64'b1001110011011110000111111101010000100100110111101010101011010110; end
            14'd13511 : begin out <= 64'b1010100110000000101001100111111110101001010111010010101111100111; end
            14'd13512 : begin out <= 64'b0010000110111111101010111011010100100100010001011010101100001110; end
            14'd13513 : begin out <= 64'b1010101011100110001010010101000000100000110000011010011110111011; end
            14'd13514 : begin out <= 64'b1010101100100000000110011101000010100000100100011010011111111110; end
            14'd13515 : begin out <= 64'b1010000111110001101010101110110100011110011111101010010110101111; end
            14'd13516 : begin out <= 64'b0010010110110010001000011111011100100100101111001010100000101001; end
            14'd13517 : begin out <= 64'b1001100010110010001010101100100000100111100100010010000011101101; end
            14'd13518 : begin out <= 64'b0010011001011010101000101110100110101010100001110001101101100011; end
            14'd13519 : begin out <= 64'b0010100101110100101001001111001010011010101010001010011000010110; end
            14'd13520 : begin out <= 64'b0010010110110101101001001000110110101011011000010010000110111000; end
            14'd13521 : begin out <= 64'b1010101011011011001001011010001100100100100010011010001011111101; end
            14'd13522 : begin out <= 64'b1010011110000000101010010000001010100011001001011001110011010110; end
            14'd13523 : begin out <= 64'b1010101110010110001010100011101010100110111011101010001101110001; end
            14'd13524 : begin out <= 64'b0010000000000110100110110110110000100100011100011010101110101010; end
            14'd13525 : begin out <= 64'b1010101110000111001010110001010100101000111110001010101100101001; end
            14'd13526 : begin out <= 64'b0001101101111000001010111001000100101000001111100010101100010111; end
            14'd13527 : begin out <= 64'b1010011010101000100111000010001010100100111011001010100110100010; end
            14'd13528 : begin out <= 64'b1010001100101011101001011111100010101011101011010010100010010100; end
            14'd13529 : begin out <= 64'b1010000010010001001010010000110010011110010111110000111101110100; end
            14'd13530 : begin out <= 64'b0010011010010011001010101110000100101001000010111010100111111100; end
            14'd13531 : begin out <= 64'b1010000100010011001000100010110110101001000111010001101000001100; end
            14'd13532 : begin out <= 64'b0010101100110010001000000011110100101010001000111001111001011101; end
            14'd13533 : begin out <= 64'b1001110001010000001010110011101000101000010111100001101110100110; end
            14'd13534 : begin out <= 64'b0010011011100001101000111110110110100000000110011010100101010100; end
            14'd13535 : begin out <= 64'b0010100100101111101001000000010110011100100110111010010110100001; end
            14'd13536 : begin out <= 64'b1010101110011000001010010111001110101011101001010010011010100111; end
            14'd13537 : begin out <= 64'b1010101110000011000011100011101010011101000111110010100100100010; end
            14'd13538 : begin out <= 64'b0010010110111010100110111001000000100100000110001001111010100111; end
            14'd13539 : begin out <= 64'b0001011010001011001010110100011010101000101001000010010001011110; end
            14'd13540 : begin out <= 64'b1001100010100100101010000101001010101001011010101001111100100110; end
            14'd13541 : begin out <= 64'b0010100010100100001001110000010110101000011101100010101111111000; end
            14'd13542 : begin out <= 64'b0010011111100010000111001110001110011111111001110010100111010110; end
            14'd13543 : begin out <= 64'b0010011001100000001010001110100010101001000101111010100010100010; end
            14'd13544 : begin out <= 64'b0010100000101101001010001101101100011110010111110010101101111101; end
            14'd13545 : begin out <= 64'b0010101110101000001001101110100000101001101000101010010001100000; end
            14'd13546 : begin out <= 64'b0010100001011101000101101001101100101000101001111010011111010000; end
            14'd13547 : begin out <= 64'b0010100001010100100111010100000010100110111111101000111011001101; end
            14'd13548 : begin out <= 64'b0010101010011100101001110101011000101000111011011010011011100100; end
            14'd13549 : begin out <= 64'b1010001100011000101010010100001010101011000011010010000101110000; end
            14'd13550 : begin out <= 64'b0010100000101011101010100010000110100111001100111010101111110001; end
            14'd13551 : begin out <= 64'b1010101100101111101010001111001000101010100100010010101101101010; end
            14'd13552 : begin out <= 64'b1010011101111001101001100001101010101000111011101010100011111010; end
            14'd13553 : begin out <= 64'b1010011000010001000110011111011010100111000000001010010001010100; end
            14'd13554 : begin out <= 64'b1010110000001000101010011111101000100101111101111010000111110000; end
            14'd13555 : begin out <= 64'b0010000010001011001010111111011010100100000010110010100011111110; end
            14'd13556 : begin out <= 64'b0010010100011110101001101110111010101011100010100010100111111101; end
            14'd13557 : begin out <= 64'b1001100001111110100111100001010110101011001011100010010010101010; end
            14'd13558 : begin out <= 64'b0010100110000011101010011100101110100000110101000010100010011011; end
            14'd13559 : begin out <= 64'b1010000011100111101010110000111010101010110000000010101100101000; end
            14'd13560 : begin out <= 64'b1010011111011000001010001101001010101010101010011010100011111000; end
            14'd13561 : begin out <= 64'b0010101000101100100100000100000110100100001110001010100111000001; end
            14'd13562 : begin out <= 64'b0010010101111011100111001110110110101001001101011001101111110011; end
            14'd13563 : begin out <= 64'b0010100000101001001010111110110000101011100011110010010100010111; end
            14'd13564 : begin out <= 64'b1001101000110111101001001010001010100011101100010010001011101000; end
            14'd13565 : begin out <= 64'b1001100110101100101010111111001010100001111011010010010111010000; end
            14'd13566 : begin out <= 64'b1010001110011111000101010010010010101010010000100010000001011001; end
            14'd13567 : begin out <= 64'b0010010011101111101010011010100110100101100111000010011100001101; end
            14'd13568 : begin out <= 64'b1010100101100101001001100000100100101000110101100010101110011011; end
            14'd13569 : begin out <= 64'b1010101110001011101010100001010100101001101001111010101101110111; end
            14'd13570 : begin out <= 64'b0010100100001101001010100011101110101010110010111010100111000111; end
            14'd13571 : begin out <= 64'b1010100100110100001010011111010000101001110101010010101111100110; end
            14'd13572 : begin out <= 64'b1010100110100111101010100001101010101011000111111010100101011110; end
            14'd13573 : begin out <= 64'b0010000100001101101010110101000100100101111110011010101011101011; end
            14'd13574 : begin out <= 64'b0010010100101100001000001011001000101010100010001010101011010101; end
            14'd13575 : begin out <= 64'b1010000011000110001001111110100010100010001000100010100100001111; end
            14'd13576 : begin out <= 64'b0010011111111111101001111101000010101010111100011001101001101010; end
            14'd13577 : begin out <= 64'b0010010110110000001001001011001010100100100011110010101001110101; end
            14'd13578 : begin out <= 64'b1010100111001001001001111110001000101010011110110010110001000000; end
            14'd13579 : begin out <= 64'b1010100000010111000111000100110100101010101110001010100011101111; end
            14'd13580 : begin out <= 64'b1010001101001010001001010001001110011110101000011010100000110110; end
            14'd13581 : begin out <= 64'b1010000110111011001001101000100100100011111111100010110000000000; end
            14'd13582 : begin out <= 64'b0010101010100001101000011010001010100101110011010010101110111010; end
            14'd13583 : begin out <= 64'b1001111001110101101000110110000000010111101100000010011010000111; end
            14'd13584 : begin out <= 64'b1010101101111110001001011100100110100110011000010010010001001001; end
            14'd13585 : begin out <= 64'b1010100100001011101010000100011100101000101001000010101011100111; end
            14'd13586 : begin out <= 64'b1010010100000101001010100010011110011100010000100010101101100110; end
            14'd13587 : begin out <= 64'b1010101111100011101010011011011100100011010110001010011011110101; end
            14'd13588 : begin out <= 64'b1010100110000001101000111011110010100100010011111010101101101010; end
            14'd13589 : begin out <= 64'b0010100011010001101010000100001010100101111011101010100110100110; end
            14'd13590 : begin out <= 64'b0010101110001000101001011010110110101010100010011010100111101101; end
            14'd13591 : begin out <= 64'b0010010011111011001000101111010000101010000101010001111111100010; end
            14'd13592 : begin out <= 64'b0010101010111110001001000010111010011110111111010001111110110011; end
            14'd13593 : begin out <= 64'b0010010011001010001010110010100110101011000101010010001001101010; end
            14'd13594 : begin out <= 64'b1010100111011011000111110010101010101000111011100010101100001010; end
            14'd13595 : begin out <= 64'b1010101011000100001001000001010110100001101011110010101000010010; end
            14'd13596 : begin out <= 64'b0010101100011010101010001011110110101000100000001010011100000110; end
            14'd13597 : begin out <= 64'b1010001000110000101010011001100100100111100000001010010011110110; end
            14'd13598 : begin out <= 64'b0010100000010010001000101101101110100110110011011010001011100100; end
            14'd13599 : begin out <= 64'b0010011011110110001010000101111110101000110011111001111000111110; end
            14'd13600 : begin out <= 64'b0010011011010001101010101001001110100110000100011010101000000001; end
            14'd13601 : begin out <= 64'b1010101100011001101010001001000110100111000101111001111110010101; end
            14'd13602 : begin out <= 64'b0010100111111101001010001000010110100100010001110010100010111111; end
            14'd13603 : begin out <= 64'b0010001011100100001010011110011000101011010011010010010010110000; end
            14'd13604 : begin out <= 64'b0010010111011010001010001010100110101001010101111010101100000011; end
            14'd13605 : begin out <= 64'b0010011001100111001010101110010110101000111001111010100000011110; end
            14'd13606 : begin out <= 64'b0010100001000111100110010000111100101010111100100010100100110110; end
            14'd13607 : begin out <= 64'b0010010001000010101000100010101100101001000101001010100110100100; end
            14'd13608 : begin out <= 64'b1001110100101101100110100111111110100111111100000001110000111011; end
            14'd13609 : begin out <= 64'b0010100000000110001010000101101100100101100001000010100001111001; end
            14'd13610 : begin out <= 64'b0010100111100001000111110010110010100000100011100010010111101111; end
            14'd13611 : begin out <= 64'b1010101000001010001010100011111100011110011000001010011001100101; end
            14'd13612 : begin out <= 64'b1010101101000011001010101111111000101000010111001001100000000110; end
            14'd13613 : begin out <= 64'b0010000001011100001010100100011110101100000000110010100101110111; end
            14'd13614 : begin out <= 64'b1010100001111000100111110000111000101011010111000001100100011001; end
            14'd13615 : begin out <= 64'b1001111110001100001010111000011100100101000001101010010010100000; end
            14'd13616 : begin out <= 64'b0010000110011010101000010000000110101001111101000010101000111011; end
            14'd13617 : begin out <= 64'b0010000101100101000111101101111110100110000110000010100110010100; end
            14'd13618 : begin out <= 64'b1010101100111001000111000111100110100100111001001010100001110110; end
            14'd13619 : begin out <= 64'b1010001101011111001000101101111000101011001110001010100110101001; end
            14'd13620 : begin out <= 64'b1010101110100110101010111101101100011101101000010001001000000001; end
            14'd13621 : begin out <= 64'b1010101111001110100111110000110000101000010110001010101011100111; end
            14'd13622 : begin out <= 64'b0010101011100101101010101001101010100111100001100010010110101011; end
            14'd13623 : begin out <= 64'b0010101011110101001000100011110000100101111100100010001110100000; end
            14'd13624 : begin out <= 64'b0010011000110010000111110101000100101100000011111010101100101100; end
            14'd13625 : begin out <= 64'b1010011000001000101001110011111100100101111110000010100001001101; end
            14'd13626 : begin out <= 64'b0010010010010010001010101101110000101011011110110010001100101001; end
            14'd13627 : begin out <= 64'b0010101011010100000111101000110100101001010001111010000001010101; end
            14'd13628 : begin out <= 64'b1010100100001010101010001011111100100101111010001010101101100001; end
            14'd13629 : begin out <= 64'b1010001001011101101010011010001010100010110000111010101111011010; end
            14'd13630 : begin out <= 64'b1010000100010001001001010001100100101010011010101010100010000110; end
            14'd13631 : begin out <= 64'b1010100010000100100111011000000100101000100011001010100001110010; end
            14'd13632 : begin out <= 64'b1010101010111010101001100010010010100011010110001001010111010010; end
            14'd13633 : begin out <= 64'b0010101101000101101010011100110010100011011101110010100001001011; end
            14'd13634 : begin out <= 64'b1001111111000101001010010101010110100100001001111010101101100111; end
            14'd13635 : begin out <= 64'b1010101010001101101000101101000110101010000010101010100000100011; end
            14'd13636 : begin out <= 64'b1010101011111110000100111000101110101001111010111010100000110111; end
            14'd13637 : begin out <= 64'b0010011000011101101001011011100000101000001100101010011000110001; end
            14'd13638 : begin out <= 64'b0001110010110000001000010000000010010110010011111010101010000001; end
            14'd13639 : begin out <= 64'b1010011100100111001010101111001110011010111001101001011111101111; end
            14'd13640 : begin out <= 64'b1010010010110010001010100100111000101011101111110010011001011110; end
            14'd13641 : begin out <= 64'b0010101111101111001010101010001000010111001000101010101011011110; end
            14'd13642 : begin out <= 64'b0010011111000001101010100001010100100000110110010010100101110100; end
            14'd13643 : begin out <= 64'b0001100110010111101000110011010010100101100011011010011010111000; end
            14'd13644 : begin out <= 64'b0010100111000111001010111001011110100111110010001010000111011010; end
            14'd13645 : begin out <= 64'b1010100100101011101010000111100110100111001010001010101000010111; end
            14'd13646 : begin out <= 64'b1010000001000000100111000000111010101000011000100010101010111000; end
            14'd13647 : begin out <= 64'b0001111100001000100011101100111110100110101011011010100011011100; end
            14'd13648 : begin out <= 64'b1010101111101110001010111011111110101001110001101010100010100000; end
            14'd13649 : begin out <= 64'b0010100001101011001010001100110000100000100010110001101110110100; end
            14'd13650 : begin out <= 64'b1010011101010101001001101110111110101011011000001010000000000010; end
            14'd13651 : begin out <= 64'b1001110110000011001010100111110000100110000010000010100000101011; end
            14'd13652 : begin out <= 64'b1010100110110101001001001000101000101001011101010010101111000011; end
            14'd13653 : begin out <= 64'b0010100101000110001010111000111100101001111010101010100111000111; end
            14'd13654 : begin out <= 64'b0010101100101011001010000000111000011110110010000010101110000011; end
            14'd13655 : begin out <= 64'b1010100001001100101010100101100010101010100110011010011101100000; end
            14'd13656 : begin out <= 64'b0010100010110011101001101101011010101010111010011010101110000101; end
            14'd13657 : begin out <= 64'b1001010111101000000010000010010110100100100011110010011101011001; end
            14'd13658 : begin out <= 64'b1010101011000001100111001001111000100000111100111010110000010000; end
            14'd13659 : begin out <= 64'b1010011111010110100110001011001000100010000100100010000011011111; end
            14'd13660 : begin out <= 64'b0010110000011110001010100000101110101010110101101010100000110000; end
            14'd13661 : begin out <= 64'b0001100111001000101001000000001100100000001011101010101001011010; end
            14'd13662 : begin out <= 64'b0010011100100111101010001010100010100100110101011010100101000100; end
            14'd13663 : begin out <= 64'b1010100001001010101001001101000000101000011000101010101001010101; end
            14'd13664 : begin out <= 64'b1010101001100110101001111010101010011100010100011010001100000110; end
            14'd13665 : begin out <= 64'b0010000111101101001010011101000110100111001110101010010001011100; end
            14'd13666 : begin out <= 64'b1010101101110101101010001011100010101000110011100010100001111010; end
            14'd13667 : begin out <= 64'b1010010001111000101001100001001110100111010111111010010011000010; end
            14'd13668 : begin out <= 64'b0010100111010101001010010000101110010100101101101010100001101001; end
            14'd13669 : begin out <= 64'b0001111000001010001001001001001110101001110010100010101100010001; end
            14'd13670 : begin out <= 64'b0001001110100011001001111111000010100110011001101010100010101000; end
            14'd13671 : begin out <= 64'b0010011000010101101010000111110000101001100101001010000000101101; end
            14'd13672 : begin out <= 64'b1010101001011001101000001100011100101010101010010001010111011010; end
            14'd13673 : begin out <= 64'b1010011011100010001001110111001100101000001100111010100111000001; end
            14'd13674 : begin out <= 64'b0001111001100001101001111000000000101001111011100010000111111000; end
            14'd13675 : begin out <= 64'b1010010101010101001010011000011100101010111110101010101011011001; end
            14'd13676 : begin out <= 64'b0010101111010101101010111101101000101001010101001010011011010000; end
            14'd13677 : begin out <= 64'b0010001010000110101010000101101000101010111101011010000110100011; end
            14'd13678 : begin out <= 64'b0010100001100100000111011000110010101010101001011010011101001010; end
            14'd13679 : begin out <= 64'b1010101010001101001001001101110100101010111001101001010000001011; end
            14'd13680 : begin out <= 64'b1010101100001100001010100110011100011110100100001010101000111001; end
            14'd13681 : begin out <= 64'b1010011111011011101010001001011110101011110010110001110011111010; end
            14'd13682 : begin out <= 64'b1010101111001101001010010100001110101011011010000001111011000111; end
            14'd13683 : begin out <= 64'b1010001111101110001010100111010010101011000011001010001110001010; end
            14'd13684 : begin out <= 64'b1010101101100010001010011100000010101010101001110010010100001101; end
            14'd13685 : begin out <= 64'b1010100100000110001001100101010010101010111010000010101010100000; end
            14'd13686 : begin out <= 64'b0010010110000110101010010001100110100101111111010010010100110101; end
            14'd13687 : begin out <= 64'b1010101011100001101010110011100000101001011100000010101100101111; end
            14'd13688 : begin out <= 64'b1010001000110010001000110000001010101001010100110010010110011000; end
            14'd13689 : begin out <= 64'b0010100001010101001001100110011100100100111111011010101101100000; end
            14'd13690 : begin out <= 64'b1010000010111110001010010110011110101011100101110010011000111001; end
            14'd13691 : begin out <= 64'b0001011111011011101010011010110110101001000001110010011001101101; end
            14'd13692 : begin out <= 64'b1001110110011011101001110010011100101011001111001010101101011001; end
            14'd13693 : begin out <= 64'b0010100110001001000110010010100000100101010111110010010100111001; end
            14'd13694 : begin out <= 64'b0010011100111100101010110100000110011110111001000010100101110001; end
            14'd13695 : begin out <= 64'b0010101000101111001000011100110100101010011100100001011010100000; end
            14'd13696 : begin out <= 64'b1010100011100010101010000101101100100111000011010001110011010111; end
            14'd13697 : begin out <= 64'b0010101000000011101000010001110010100111111101111010010010010011; end
            14'd13698 : begin out <= 64'b1010100010010100101010000011001110011001010011001010001110001100; end
            14'd13699 : begin out <= 64'b1010100100000111001010010010110010100110001100011010101100001011; end
            14'd13700 : begin out <= 64'b0010010010100011100111100111111010101000000101011010101111010001; end
            14'd13701 : begin out <= 64'b1001110000011111001001010000100010101001011011100010001101101011; end
            14'd13702 : begin out <= 64'b1010011001000100101001001001110100101100010000110010011011001011; end
            14'd13703 : begin out <= 64'b0010010000101100001001000100111000011001111111001010101010110100; end
            14'd13704 : begin out <= 64'b1010101101011111101001011111111000101010000111111010100011110101; end
            14'd13705 : begin out <= 64'b1010010000110100001011000101001000101001001010101010000101010110; end
            14'd13706 : begin out <= 64'b1010101010011110101010000110011100011111011001001010101111100101; end
            14'd13707 : begin out <= 64'b0010100100011100101001011100101000101010011110000010101011111111; end
            14'd13708 : begin out <= 64'b0010011100111110001000010010110100100010001001100010100111100001; end
            14'd13709 : begin out <= 64'b0001100100001000101010011000110100100100100001101010011110010100; end
            14'd13710 : begin out <= 64'b1010100100000010101010111100111000011000011101100010101011001110; end
            14'd13711 : begin out <= 64'b0010101010001110101010111110010000101011101000011001101111001000; end
            14'd13712 : begin out <= 64'b0010011000101001001000011111010110011111011110111010101010010000; end
            14'd13713 : begin out <= 64'b0001001001011010101010100101001000101010001111110010010000111010; end
            14'd13714 : begin out <= 64'b0010101111110100001001101001101010100110111001110010011001000100; end
            14'd13715 : begin out <= 64'b0010100000010101101010101100011110100111100111111010110000011010; end
            14'd13716 : begin out <= 64'b1010101101001010101010010100111100101011101100101010101100101110; end
            14'd13717 : begin out <= 64'b0010000110001101100011100000000100101010010010011001110011110100; end
            14'd13718 : begin out <= 64'b1010010001101010001000000111010110100110001111111010101000001011; end
            14'd13719 : begin out <= 64'b0010101000000000101001110111000100101001011000100010000111000110; end
            14'd13720 : begin out <= 64'b0010000101010011001000011111010000010101111000111010101010000000; end
            14'd13721 : begin out <= 64'b0010011101111100001001111011110100100111001111110010000110000101; end
            14'd13722 : begin out <= 64'b0010100011011111001010001101111100100000010001011010100100001010; end
            14'd13723 : begin out <= 64'b1010100011110000101000010101110100101001000100100000110111011000; end
            14'd13724 : begin out <= 64'b0010101011010000100110101111101110101100010011000010101101001101; end
            14'd13725 : begin out <= 64'b1010000010101010100101101100011100100101110001101010100110101001; end
            14'd13726 : begin out <= 64'b0010011100110101001000001000001010101000011011000010110000001011; end
            14'd13727 : begin out <= 64'b0001110010010001100101111110100000011111111111101010011001111000; end
            14'd13728 : begin out <= 64'b0001110100110101001010000110001010100111101011011010101111011100; end
            14'd13729 : begin out <= 64'b1001110010101001001010010100110010101000011101010010101110001001; end
            14'd13730 : begin out <= 64'b0010100111101111101010110011101100100011011000010010010111110110; end
            14'd13731 : begin out <= 64'b1010101001010011101001010101000010101100001101100010011100110001; end
            14'd13732 : begin out <= 64'b1010010100101111001010001101011100101010000011100010100101011000; end
            14'd13733 : begin out <= 64'b1010010101100100001010100111010000101010100100001010010011100001; end
            14'd13734 : begin out <= 64'b1010101110000001001001011011110100100001101011110010101001101001; end
            14'd13735 : begin out <= 64'b1010011101111101001010001111101010101001100110100010101101011011; end
            14'd13736 : begin out <= 64'b0010101010101010001001000000111010100101000110111010000101010100; end
            14'd13737 : begin out <= 64'b1010101000010101001010000100001000101001000010111010010111010110; end
            14'd13738 : begin out <= 64'b1010001111000011001001001000101100101000011010110010010110000101; end
            14'd13739 : begin out <= 64'b1010010010100100001001111000010010101001000001001010101101110101; end
            14'd13740 : begin out <= 64'b1010010110000001101010111110011000101001101101111010100111101100; end
            14'd13741 : begin out <= 64'b0010011101100011101000100011101100101010111000000010100000100001; end
            14'd13742 : begin out <= 64'b1010100000001000000111100000101100101010010110110010110000011101; end
            14'd13743 : begin out <= 64'b0010011000011011001010100110110010011000110001110010001011110000; end
            14'd13744 : begin out <= 64'b0010011011111110001001100000110010100111001010100010011010101110; end
            14'd13745 : begin out <= 64'b0010010111000000001010000001101100100101110011010010010111101001; end
            14'd13746 : begin out <= 64'b1010011011010101100111000010001110100110111000110010000101101100; end
            14'd13747 : begin out <= 64'b0001110110101011001001011101011100100100101101100010010111010011; end
            14'd13748 : begin out <= 64'b1010100110010101001001011011011010101001111100110010001010100110; end
            14'd13749 : begin out <= 64'b0010100010010011100101010001101000011110000111101010100111001111; end
            14'd13750 : begin out <= 64'b0010011011111100101010001010110010101011011101110001111111011001; end
            14'd13751 : begin out <= 64'b0010101000010100101010010101000110100101000001100010011010001111; end
            14'd13752 : begin out <= 64'b0010100111010100100110001110000000100110001000110010100010010100; end
            14'd13753 : begin out <= 64'b1010100110010101001010110100101100011100110011111010100000111101; end
            14'd13754 : begin out <= 64'b0001110110011000001010000011101000101000000011101010101111001110; end
            14'd13755 : begin out <= 64'b1010100000010110100101010101100010011010010001010010110001001110; end
            14'd13756 : begin out <= 64'b1010011011010110101010011111100110100001001101010010011111111101; end
            14'd13757 : begin out <= 64'b0010011010011001101001010001101010100110101100001010001000000010; end
            14'd13758 : begin out <= 64'b1010100011001111101000111110011100100101001111101010100111100110; end
            14'd13759 : begin out <= 64'b0010000111010111101000001000110010101010011000101010010010011000; end
            14'd13760 : begin out <= 64'b0010100111001000001001110110100110101001000101110010000101010110; end
            14'd13761 : begin out <= 64'b0010101110001100101010011111001110101001000000011010001010010100; end
            14'd13762 : begin out <= 64'b0010011000001010101010111101111000100101111000011010100000110110; end
            14'd13763 : begin out <= 64'b1010101100001100100111010000011110100001101110000010000100010000; end
            14'd13764 : begin out <= 64'b1010010100101000101001001101000000101001000101111010011010011011; end
            14'd13765 : begin out <= 64'b0010101010100010001010000110010010101001101111101010100100110100; end
            14'd13766 : begin out <= 64'b0010101000011001101010010101000110011110001010110001111110101101; end
            14'd13767 : begin out <= 64'b1010000010011011001001110101111000100101110101110010101011101111; end
            14'd13768 : begin out <= 64'b1001110100111101101010010010100010100110101101000010100010111111; end
            14'd13769 : begin out <= 64'b0010011110101111001000101001011100100100110101101010100010111010; end
            14'd13770 : begin out <= 64'b0010001010001000101010011101101010101011000000110001100100101010; end
            14'd13771 : begin out <= 64'b1010011010000000001001011111011000101001101000010010100000001110; end
            14'd13772 : begin out <= 64'b1010100001100111001000000001100100101001000010100010100110110110; end
            14'd13773 : begin out <= 64'b0010101110000101101001000100001000101000101001000010001010010000; end
            14'd13774 : begin out <= 64'b0010101101010110001001110111110110101000111001110010100100111110; end
            14'd13775 : begin out <= 64'b0010010111111111101001011011110100101011011100110001110011011110; end
            14'd13776 : begin out <= 64'b1001110011111110001010100001011000010100011110011010101110100100; end
            14'd13777 : begin out <= 64'b0010010011101011101010110110110010100111101011111010000001001001; end
            14'd13778 : begin out <= 64'b1010101100011011101001101011101100100101001001010010010110001011; end
            14'd13779 : begin out <= 64'b0010101100001011001001000000001100101000010000000010100010100101; end
            14'd13780 : begin out <= 64'b1010101000010110101010001000111100101001110100001010101001111100; end
            14'd13781 : begin out <= 64'b1001110010010101101001000001010000100100101111111001100001001001; end
            14'd13782 : begin out <= 64'b1010101001000011001010010001110000100100110101111001101100001011; end
            14'd13783 : begin out <= 64'b0010011000010100101010001101110100101001001100000010000101010110; end
            14'd13784 : begin out <= 64'b1010000101001111101000101101111100100001000111110010010010000110; end
            14'd13785 : begin out <= 64'b0010000111101000101001100000110110100110010100110010100011110000; end
            14'd13786 : begin out <= 64'b1010101001011001101000110100011100011100010011011010100100111101; end
            14'd13787 : begin out <= 64'b0010101000110000101010000001110000101010110100110010100101010110; end
            14'd13788 : begin out <= 64'b1010010010111101001001011111110010100101011011011010011100101011; end
            14'd13789 : begin out <= 64'b0010101111110100101000001110101100100101110000010001110101011111; end
            14'd13790 : begin out <= 64'b0010101000111010001010101111011100101010110001011010011001001000; end
            14'd13791 : begin out <= 64'b0001010011110000001010110001100010101000000001000010100111011010; end
            14'd13792 : begin out <= 64'b1010100000110100001001100010001110101000101110010010101000001101; end
            14'd13793 : begin out <= 64'b0010101010000111001000001111011100100011110000110010011111011110; end
            14'd13794 : begin out <= 64'b1010001100110011001010011001110000011110110001101010101101110111; end
            14'd13795 : begin out <= 64'b0010100010111100101010101111100010100110001110011010100100011010; end
            14'd13796 : begin out <= 64'b1010100111010001001001101111101110100111000111000010010001011011; end
            14'd13797 : begin out <= 64'b1010101010010010001010100101110110100101111001000010011000110101; end
            14'd13798 : begin out <= 64'b1010010001000100101000001100011110100101001111000010101000001001; end
            14'd13799 : begin out <= 64'b0010000111000001101010100100001110101001010000100010101111100111; end
            14'd13800 : begin out <= 64'b1010101010011111100101011100001000100101100110101010101010010101; end
            14'd13801 : begin out <= 64'b1010001011110011101000001100111010100101001100100010000100001100; end
            14'd13802 : begin out <= 64'b1010100101101010101010000000000100101010111010000010001011110100; end
            14'd13803 : begin out <= 64'b0010010011011111001010001000010010100111001110000010110000000010; end
            14'd13804 : begin out <= 64'b1010101001101011101010100100101010101010100111110010100111101011; end
            14'd13805 : begin out <= 64'b1010101111000011001000001100001100100010000000011010101000101101; end
            14'd13806 : begin out <= 64'b1010100001000100101000101110011000001100000100100001101110101001; end
            14'd13807 : begin out <= 64'b0010100001010110001000100001101110101010101110110010100010011010; end
            14'd13808 : begin out <= 64'b0010101101110110001000011000111010101010011111011010000111001010; end
            14'd13809 : begin out <= 64'b0010000010101110001010001000000010011110100100010010100101101010; end
            14'd13810 : begin out <= 64'b1010010001000101001010001011000000101011000110101010011110011110; end
            14'd13811 : begin out <= 64'b0001101111101010001010000001111000101010100011111010101010011010; end
            14'd13812 : begin out <= 64'b0010100111011000101010110010011110100100101111110001011110100010; end
            14'd13813 : begin out <= 64'b0010100110010101001010011100100100011110101110100010110000111110; end
            14'd13814 : begin out <= 64'b0010010101101010101010110101010110100001101000100001111101001100; end
            14'd13815 : begin out <= 64'b1010000110100111000111111101110010101000000000101010010101000110; end
            14'd13816 : begin out <= 64'b1010100101000010001010011000000100101000100000100010001100110111; end
            14'd13817 : begin out <= 64'b0010011011010111101011000000111000011110100010000001110011010100; end
            14'd13818 : begin out <= 64'b0010100011111000101010011001100110100101010110111010000100111011; end
            14'd13819 : begin out <= 64'b1001111110100011101010011001010100100100000001110010100110101011; end
            14'd13820 : begin out <= 64'b1010101001001001000110011101101010101000110100011010101101011101; end
            14'd13821 : begin out <= 64'b1010011001100111000111001010000100101001111110011010100010100111; end
            14'd13822 : begin out <= 64'b1010101110101010001010111001110010100010100100011010101000000011; end
            14'd13823 : begin out <= 64'b1010000110111101001010010011001010100010111100100010110000111111; end
            14'd13824 : begin out <= 64'b0010000111011101101010110000000110100111110110110010011101110111; end
            14'd13825 : begin out <= 64'b1010101101000010101000100010100100101011100010011010000001111011; end
            14'd13826 : begin out <= 64'b0010101011001101001000000000101100100000011001111010101101110101; end
            14'd13827 : begin out <= 64'b0010101100011110001010011000100010100000111000100010101100011111; end
            14'd13828 : begin out <= 64'b0010001110111010001001100111010010100001011011001010100000001001; end
            14'd13829 : begin out <= 64'b0001111111011001101010001000001000011110101110101010010101110001; end
            14'd13830 : begin out <= 64'b1001001010100000101010011111000000101011001111011010011011011001; end
            14'd13831 : begin out <= 64'b0010100100100100001010000000000100101011000011010001111010011001; end
            14'd13832 : begin out <= 64'b0010100111001111001001000111110010101010111000101001100100000000; end
            14'd13833 : begin out <= 64'b0010011101001101001010100101101000100111000100101010101011110011; end
            14'd13834 : begin out <= 64'b0010010110000000000110001000100000011000111111011010110000011000; end
            14'd13835 : begin out <= 64'b0010101111110100001001011011001000011010010000011010100110101100; end
            14'd13836 : begin out <= 64'b0010011001011110101010001110011110011101110111010010010111000000; end
            14'd13837 : begin out <= 64'b0010101110000111101010001011011100100110111111111010101000100011; end
            14'd13838 : begin out <= 64'b0010100010101000101010110101111010100001000111010010100011010010; end
            14'd13839 : begin out <= 64'b1010001000010010101010011101100100100110000011100010011101110011; end
            14'd13840 : begin out <= 64'b0010101011110111101000000001100010101010000111110010011101011001; end
            14'd13841 : begin out <= 64'b1010011111100111101001101001100010010010100111000010100001111111; end
            14'd13842 : begin out <= 64'b1001010010010101001001110010011100011100111000000010101011001111; end
            14'd13843 : begin out <= 64'b1010000010110010101010101101101110100101001110011010101111110000; end
            14'd13844 : begin out <= 64'b1010101110110110001010100001111010100001100010011010101010001110; end
            14'd13845 : begin out <= 64'b1010100111000011101010000110011000100011011100100010100110101001; end
            14'd13846 : begin out <= 64'b1010010100010100001001101010011110010101010101000001111010000111; end
            14'd13847 : begin out <= 64'b1010100010000001001010101100110110101010010001001010101100101011; end
            14'd13848 : begin out <= 64'b0010101000100110101001101100011100101001001011101010101011110001; end
            14'd13849 : begin out <= 64'b0010010001111110001010000001000010101010111101111001101011001101; end
            14'd13850 : begin out <= 64'b1010100111101001101010011101011100101010100100011010100011010011; end
            14'd13851 : begin out <= 64'b1010010101010101001010110000001100100111011010110010010001110000; end
            14'd13852 : begin out <= 64'b1001101111101010101001101010000010100011101101000001111000110001; end
            14'd13853 : begin out <= 64'b1010101000111111001010011110101110101000110000001010100100000101; end
            14'd13854 : begin out <= 64'b0010101011010111001001010111010000101000001111001010101100110011; end
            14'd13855 : begin out <= 64'b1001000110111011001001010000101100101001001110101010100001101101; end
            14'd13856 : begin out <= 64'b1010100110001000001010100101110100101011011010101010101010110100; end
            14'd13857 : begin out <= 64'b1010100110110111000110001101100100100100001110111010011001000010; end
            14'd13858 : begin out <= 64'b1010001011111010001000010101010100100110001010011010010101001010; end
            14'd13859 : begin out <= 64'b0010101110101010101010100010001010101010000010101010101101100011; end
            14'd13860 : begin out <= 64'b1010101001010100101010111001111010101011110101001010100001110111; end
            14'd13861 : begin out <= 64'b0010001101101010101001101010010100101011100111101010110000001110; end
            14'd13862 : begin out <= 64'b0001110111101110001001010110101110101001110000001001000001011001; end
            14'd13863 : begin out <= 64'b1010011110011001101010000000101100100111001011110010010101101100; end
            14'd13864 : begin out <= 64'b0010010011011111101001111111010100101010000011111010101100101111; end
            14'd13865 : begin out <= 64'b1010010100001000001000000111001000011111101000011010100110101100; end
            14'd13866 : begin out <= 64'b1010100011000111101010010000100100101011110111110010101011001000; end
            14'd13867 : begin out <= 64'b0010010101000110001000100111011100101011100111111010000011000010; end
            14'd13868 : begin out <= 64'b0010001011011100101010101010010100101011110011001010001001111011; end
            14'd13869 : begin out <= 64'b1010101011001011101001011010100000011001010010010010011111001001; end
            14'd13870 : begin out <= 64'b0010110000000111001000001101110000101011010111011010100110000100; end
            14'd13871 : begin out <= 64'b1010001000110011001001101100001100101011001101110010100110011001; end
            14'd13872 : begin out <= 64'b1010000111100011101000001101110010101000000101110010101110000111; end
            14'd13873 : begin out <= 64'b1010101010011101101010111000111010101000111100010010010011011010; end
            14'd13874 : begin out <= 64'b1010001011011000101010000000100000100101000111011010000000111110; end
            14'd13875 : begin out <= 64'b0010100001110010001010110101110110100101101010111010101010101110; end
            14'd13876 : begin out <= 64'b0010100101100110001010110010010100100111010100010010100001011001; end
            14'd13877 : begin out <= 64'b0010100011111001101001101001100110101010101111100010101100100110; end
            14'd13878 : begin out <= 64'b1010011000110001001000100001001010011101000001110010011111010011; end
            14'd13879 : begin out <= 64'b1010010010101011101010101010100000001001110010000010100101111111; end
            14'd13880 : begin out <= 64'b0010101100010011101000111110100000100001011110001010100111100010; end
            14'd13881 : begin out <= 64'b1001011001000010101010100110010110101000111000101010101110000001; end
            14'd13882 : begin out <= 64'b1010101101011110101001000001010110101011010111100010000011110011; end
            14'd13883 : begin out <= 64'b1010100110101110001001011111111000101000111110000010101001111110; end
            14'd13884 : begin out <= 64'b0010100110001100001001010111011010101010001100101010101111111011; end
            14'd13885 : begin out <= 64'b0010101111100110100101110100011000101001000011000001101000101001; end
            14'd13886 : begin out <= 64'b1010011101100011001010010111101000101011010011100001000010010101; end
            14'd13887 : begin out <= 64'b0001000111110111101010011010100100101010001100101010011001011111; end
            14'd13888 : begin out <= 64'b1010011100111000001001100111000110100101000011111010100010000001; end
            14'd13889 : begin out <= 64'b0001011011011010000110100001001010011110011011111010100100110110; end
            14'd13890 : begin out <= 64'b1010000100010110101010111111011010011101100111011010011000000011; end
            14'd13891 : begin out <= 64'b1010101011010111000111011100011110011001100001000001101010010010; end
            14'd13892 : begin out <= 64'b0010100011101011001010111110011110101000001110011010101001101101; end
            14'd13893 : begin out <= 64'b1001110000110001001001010011000010101010011000101010101000100101; end
            14'd13894 : begin out <= 64'b0001101011011111001010000111101110101011110000011010011101010100; end
            14'd13895 : begin out <= 64'b1001100010011000101010101011110000100101111101000010101011101100; end
            14'd13896 : begin out <= 64'b1010101010110001101010110010010100100101010101100010100010101110; end
            14'd13897 : begin out <= 64'b1001111010100100001001101001111100101000001101101001111010001111; end
            14'd13898 : begin out <= 64'b1010001100010110101001001000101010100100011101011010101111011100; end
            14'd13899 : begin out <= 64'b0010100011110010001000111100101010100011101011001001111110010011; end
            14'd13900 : begin out <= 64'b0010011001111110001010100101000000100001100100111010001100101010; end
            14'd13901 : begin out <= 64'b1010011101101110001010010101001100101001000111100010100100000010; end
            14'd13902 : begin out <= 64'b0010010011100011001001111001000100100010100111001010100000011100; end
            14'd13903 : begin out <= 64'b1010010011110011001010001100110010101000101000100010010011010100; end
            14'd13904 : begin out <= 64'b0010100100101001001010111011011010101010100101001010100100001011; end
            14'd13905 : begin out <= 64'b0010100011110000101010001000111110101000101000111010001110010111; end
            14'd13906 : begin out <= 64'b1010100110010001101010010111010110011110101011001010100000110111; end
            14'd13907 : begin out <= 64'b1010110000110110101010100101110100101000011011101010001110101100; end
            14'd13908 : begin out <= 64'b0010101001011101001010001011001100011010110000011010101111101001; end
            14'd13909 : begin out <= 64'b1010101100111100001010101010001010101011111111111001011001101111; end
            14'd13910 : begin out <= 64'b0010001000011001001000001100010000011010100111010010001001000000; end
            14'd13911 : begin out <= 64'b0010101101010011001010010100111010101010101110010010010110110001; end
            14'd13912 : begin out <= 64'b1010010110101011101001000110100100101001111010000010100111011100; end
            14'd13913 : begin out <= 64'b0001110001111000001000010001100110011011101011100010101011111001; end
            14'd13914 : begin out <= 64'b0010001100111010100111110000010110100100011001011001110110101011; end
            14'd13915 : begin out <= 64'b0010100111101011101010100101000000101001010110001010100011110101; end
            14'd13916 : begin out <= 64'b0010011011001001101010010101101010101000000010101010100000000111; end
            14'd13917 : begin out <= 64'b0010010011101100101010011101011000011010010010000010101101010010; end
            14'd13918 : begin out <= 64'b1010100111101001001010000001100100011110111101000010000000011111; end
            14'd13919 : begin out <= 64'b1010110001110010101000001100000010101000110010101010011011001001; end
            14'd13920 : begin out <= 64'b1010010010011010001010100111100010100101010001111010100110111001; end
            14'd13921 : begin out <= 64'b0010011011111101101010011101111000100111100110010010010011000010; end
            14'd13922 : begin out <= 64'b0010100101100001001000000101110010101001110001001010001111100100; end
            14'd13923 : begin out <= 64'b0010011111111111101010110000111010101000001001001010100100101101; end
            14'd13924 : begin out <= 64'b1010010000011111001010000100110000101001100010001010011000000100; end
            14'd13925 : begin out <= 64'b0010101011011111001010101101110110101000110110001010101101011110; end
            14'd13926 : begin out <= 64'b0010010010101111000111111110010000100110010000101010100101111011; end
            14'd13927 : begin out <= 64'b1010101011100111001000010000000110101010010111111010101111010000; end
            14'd13928 : begin out <= 64'b1000000001110111001000001001000010101011101001010010101011011001; end
            14'd13929 : begin out <= 64'b1001110000101111101010010001111100100011000110100010001000100000; end
            14'd13930 : begin out <= 64'b0010000000100010001010010001001000101011111111101010100011110111; end
            14'd13931 : begin out <= 64'b0010101001110110001010100011110100101001011100101010101111000110; end
            14'd13932 : begin out <= 64'b0010001000001010001010111000111010100111111001110010001110100101; end
            14'd13933 : begin out <= 64'b0010000010100100001001101101001010101011010111001010100011001100; end
            14'd13934 : begin out <= 64'b1010101001111010101010110001010110100011001110101010100001110100; end
            14'd13935 : begin out <= 64'b0010010011101111101010000010110010100000011111110001000100011111; end
            14'd13936 : begin out <= 64'b0001011001110011101000011001000000101000110011100010101011011001; end
            14'd13937 : begin out <= 64'b0010101010111011101001011100011010100110110011001010101010010111; end
            14'd13938 : begin out <= 64'b0010001111111101100111100111111010100100011111100010101111010111; end
            14'd13939 : begin out <= 64'b0010100001010011001010111001010010100110101111100010010110000001; end
            14'd13940 : begin out <= 64'b1010100101010101101001001111011010010000100011001010000111001111; end
            14'd13941 : begin out <= 64'b1010101000011010101001101110111100101010000000110010100101000000; end
            14'd13942 : begin out <= 64'b0010010111000010001010011100100000100101101001000010000111111111; end
            14'd13943 : begin out <= 64'b0010100111110010001001100110111000101010111110000010101000001110; end
            14'd13944 : begin out <= 64'b1010000110100100100110111011100000100001000100010010100001100000; end
            14'd13945 : begin out <= 64'b0010101100101011101001010000110000101000011000010010010101110110; end
            14'd13946 : begin out <= 64'b0010011011000011101001101010000110101011000010010010101010101110; end
            14'd13947 : begin out <= 64'b1010100110001110001010001101010000101001001111001010100010011001; end
            14'd13948 : begin out <= 64'b1010101110100101001010111110111010101011101001000001110100101001; end
            14'd13949 : begin out <= 64'b1010101001110011101010011000110000011111010110000010100000010011; end
            14'd13950 : begin out <= 64'b0010100100010110001000111100010100011110011101101010001011000101; end
            14'd13951 : begin out <= 64'b0010100111100011001010111110000100100101111111011010010110010111; end
            14'd13952 : begin out <= 64'b0010100011001100001010011100110000101010100111001010100100000010; end
            14'd13953 : begin out <= 64'b1010100011011011001010100001100000100110100110001010101101111000; end
            14'd13954 : begin out <= 64'b0010010001100100001001100001011100101010111001101010101011010100; end
            14'd13955 : begin out <= 64'b0010011100100000001000010000001000100111011000110010100011010010; end
            14'd13956 : begin out <= 64'b1010011110110101001010111010010010011101010110101010011010100000; end
            14'd13957 : begin out <= 64'b1010000011101011101010100011010110101001110010101010100101011001; end
            14'd13958 : begin out <= 64'b1010101000100000001010000001001100100100101100000010010110111111; end
            14'd13959 : begin out <= 64'b0010101010010111101010010011010000101000101110001010100100001010; end
            14'd13960 : begin out <= 64'b1010000101100001101000000110110100101001111110101010100010010110; end
            14'd13961 : begin out <= 64'b1010000010000010001010100000110100101000111100001010010010000101; end
            14'd13962 : begin out <= 64'b1001101111110010101000010011010110101011011000001010100010010111; end
            14'd13963 : begin out <= 64'b0001110010110010100110000001011000100100110110010010100000001010; end
            14'd13964 : begin out <= 64'b0010100011011101001001011110100000101000011000100010001001101001; end
            14'd13965 : begin out <= 64'b1010101101001110101001011011110000100101100000011010000011100101; end
            14'd13966 : begin out <= 64'b1010000100100110101010111100101100011100010101110010010000100110; end
            14'd13967 : begin out <= 64'b0010101011110000101001100011001100100100010101100010011101110110; end
            14'd13968 : begin out <= 64'b1010010011011101001010011100111000100111010110101010010000010000; end
            14'd13969 : begin out <= 64'b1010010101001110001010111111101010011110010101110001011010110101; end
            14'd13970 : begin out <= 64'b0010011101110000101010011001111010101001100101011010101001011000; end
            14'd13971 : begin out <= 64'b1010100100111000001010111001110010100100110011110010101011100101; end
            14'd13972 : begin out <= 64'b0010101010010001101010101010100000101010100001100010100111111001; end
            14'd13973 : begin out <= 64'b1010101110101110000111010100110010100000010101010010001011001101; end
            14'd13974 : begin out <= 64'b1001110001101001100111101111000010101010000101010010101010101000; end
            14'd13975 : begin out <= 64'b1010100101101011001010100101011000100011111100111010101101101001; end
            14'd13976 : begin out <= 64'b0010101100110010101010010110101100011111001010110010100001100011; end
            14'd13977 : begin out <= 64'b0010100101101110101010000000111010010110000110100010100010001111; end
            14'd13978 : begin out <= 64'b1010101001000110101001111011100010100111001000111010010110001100; end
            14'd13979 : begin out <= 64'b0010010110000101101010001001001100101010000110101010101101000001; end
            14'd13980 : begin out <= 64'b1010101000110010001010000001000110011011001010000010101111110001; end
            14'd13981 : begin out <= 64'b1010001001000100101010010100001000100110111001111010101010001111; end
            14'd13982 : begin out <= 64'b0010000101011101101010100111001010100001010001110010101110011101; end
            14'd13983 : begin out <= 64'b1001111000000101101001001100001110100010001011010001110010101101; end
            14'd13984 : begin out <= 64'b1010101110101011001001010000101000101000101000110010010011100100; end
            14'd13985 : begin out <= 64'b0001110111011110000111101111010110100010101001111010100010100110; end
            14'd13986 : begin out <= 64'b0010101111100011001010001011011100101000111010110010011011010010; end
            14'd13987 : begin out <= 64'b0010001100000000101001111001101010101001000111100010010101001101; end
            14'd13988 : begin out <= 64'b1010010010011101101010111000101100101010101010000010101010011010; end
            14'd13989 : begin out <= 64'b0010010000110011000111101011011100101010011111100010101001111110; end
            14'd13990 : begin out <= 64'b0010101110011000001010101010001000101000000000100001000101111000; end
            14'd13991 : begin out <= 64'b1001111100111100001001101010100000100110101110011010011001000110; end
            14'd13992 : begin out <= 64'b0010100100010101001010111111111000100000100101101010100110011101; end
            14'd13993 : begin out <= 64'b0010011011110010101000100100000000101000010010001010001000100000; end
            14'd13994 : begin out <= 64'b1010010010010011001000111010001100101010010100001010010110110010; end
            14'd13995 : begin out <= 64'b0010001001001011101001001110010100101000110001100010011001001110; end
            14'd13996 : begin out <= 64'b0010101001101100001001111011111000101000000100110010010101100010; end
            14'd13997 : begin out <= 64'b0010101000111001101010101100010100100010101010000001001010111100; end
            14'd13998 : begin out <= 64'b1010100111000011101010111011101100100101101111111010100110011111; end
            14'd13999 : begin out <= 64'b1010101111111100000101011110111010101011010011011001111000011011; end
            14'd14000 : begin out <= 64'b1010010000111010101001100001000100101001010101011010000101011111; end
            14'd14001 : begin out <= 64'b1010011110010101001001100111111110101000000110001010001110010111; end
            14'd14002 : begin out <= 64'b1010101001101000101001011101101010101010010101011010101000011001; end
            14'd14003 : begin out <= 64'b0010011010101010001001110000001000100001011100100010100111010111; end
            14'd14004 : begin out <= 64'b1010010111001001101000111000111010101010010000011010101101101111; end
            14'd14005 : begin out <= 64'b1010011000001001001010101111000010100101101010001010101011101001; end
            14'd14006 : begin out <= 64'b1010101110000000101010101110011000100100110101100010100111111011; end
            14'd14007 : begin out <= 64'b0010100111100111001010110010100000101011101101001010010110000000; end
            14'd14008 : begin out <= 64'b1001110011111010101001111110101110100000011001001010010001001100; end
            14'd14009 : begin out <= 64'b1010101100101100001010010000010110011110001000111010001110110010; end
            14'd14010 : begin out <= 64'b1010010010110010001001011111110000100000001101111010000110001101; end
            14'd14011 : begin out <= 64'b1010001101111101101010100000110000011111000110011010010011111010; end
            14'd14012 : begin out <= 64'b0001111011101100100101000010101000101001000111110010101100101110; end
            14'd14013 : begin out <= 64'b1001100100000110001010110011110100101000111110000010000111111000; end
            14'd14014 : begin out <= 64'b0010001001110001001010100011000100101011110000111010010001011000; end
            14'd14015 : begin out <= 64'b1010100010011110101010010000001000101010100111001001111001101000; end
            14'd14016 : begin out <= 64'b0010011010111110001001100000010000010100000000011000101111100000; end
            14'd14017 : begin out <= 64'b1010011101001101101010101110001100100110011011011010100001111000; end
            14'd14018 : begin out <= 64'b0010011101001000101001010100010110101000101001110010100000100100; end
            14'd14019 : begin out <= 64'b1010000101110111001001101010010010101011100001100010100010001011; end
            14'd14020 : begin out <= 64'b0010001011001010001010111011111000100101100110100010100111010010; end
            14'd14021 : begin out <= 64'b1010100010000101001010000011011110010111101011110010011000011001; end
            14'd14022 : begin out <= 64'b0000101101000100001001000101101000100111100100000010101011010111; end
            14'd14023 : begin out <= 64'b0010010110101111001001100110110010101000100010100001011001101100; end
            14'd14024 : begin out <= 64'b0010000111100000101010011101010000100010001110011001110110011100; end
            14'd14025 : begin out <= 64'b1010101101000110001000011101001010101001001000000010101101100101; end
            14'd14026 : begin out <= 64'b0010000110111110100111110101101110100111101110110010010010111111; end
            14'd14027 : begin out <= 64'b1001111000001101001000010111110100100011111111000010011101101111; end
            14'd14028 : begin out <= 64'b0010101011000011001010110000101100100000100011000010101111011100; end
            14'd14029 : begin out <= 64'b0010100110011101001001011000001010101010010001110010011011100101; end
            14'd14030 : begin out <= 64'b1010011011110101101001010110001010100110101000111010100111010001; end
            14'd14031 : begin out <= 64'b0010011100000110101010000110101100101001100111000010101001111011; end
            14'd14032 : begin out <= 64'b1001101010110000101000011000110000100100100110010010100111011001; end
            14'd14033 : begin out <= 64'b1010000101000000101010101101111110100100101001001001001100001111; end
            14'd14034 : begin out <= 64'b1010000101101000101010010110011100011110111000000010000111001101; end
            14'd14035 : begin out <= 64'b1010100011000111101001110001100110101011010100010001101101111100; end
            14'd14036 : begin out <= 64'b1010101011001001101001000101101010011101001100001001111101011001; end
            14'd14037 : begin out <= 64'b0010101101101001101010001100101100011111010100000010000001111100; end
            14'd14038 : begin out <= 64'b1010100011011100001001000101001100101000001010110000011110000110; end
            14'd14039 : begin out <= 64'b1010000101010111001000101011001000101010111111001010011001100110; end
            14'd14040 : begin out <= 64'b1010100110010010101010111100011000011110100011010010100110000100; end
            14'd14041 : begin out <= 64'b1010101001001011101001000001011000101001100111111010101001011111; end
            14'd14042 : begin out <= 64'b0010101111011011101010110000000000100011101001101010101011110001; end
            14'd14043 : begin out <= 64'b0010100100101011001000100001001110101010110011111010011000011101; end
            14'd14044 : begin out <= 64'b0010100000100111001010010110100100100001010000011010001011001011; end
            14'd14045 : begin out <= 64'b1010010101011000001010001000111110100010100110010000110100111000; end
            14'd14046 : begin out <= 64'b0010101010101111101010001101001110011001100000111010101111100101; end
            14'd14047 : begin out <= 64'b1010110000011110101010111111111110011100000110001010001011100100; end
            14'd14048 : begin out <= 64'b0010000100001110100111110110000110101000000001110010001100111000; end
            14'd14049 : begin out <= 64'b0010011011001101001001010011000010101011101000011010101010101110; end
            14'd14050 : begin out <= 64'b0010100100100101101010010110010000100100010011111010000000101011; end
            14'd14051 : begin out <= 64'b1010100101010110101010111001010010101001010101101010101000101001; end
            14'd14052 : begin out <= 64'b0010000111000000101010101101010010100011011110000010001001011000; end
            14'd14053 : begin out <= 64'b0010100010011011001010010000101110100111100100111010001100100010; end
            14'd14054 : begin out <= 64'b1010100100101011100110011001001000100101101111110010100110100011; end
            14'd14055 : begin out <= 64'b1010101000011001101001010111110100101000011111000010011011010001; end
            14'd14056 : begin out <= 64'b1010001001011101101010010110111100101001000010010010010000100100; end
            14'd14057 : begin out <= 64'b1010011111101111101010000010010110011100101001010010010101110101; end
            14'd14058 : begin out <= 64'b1010001100101111101010001000100100100010000011111010011100011000; end
            14'd14059 : begin out <= 64'b1010100001011111101010000101011110100101000011100010100111101010; end
            14'd14060 : begin out <= 64'b0001010111100000001001000101000010011010010011111010100000101001; end
            14'd14061 : begin out <= 64'b1001101101011100000111110101000000010100011101010010010101000111; end
            14'd14062 : begin out <= 64'b1010101101111100001010000001110100100110110110110010100011110101; end
            14'd14063 : begin out <= 64'b0010011000100011101010001110100100100010101001001010101111011100; end
            14'd14064 : begin out <= 64'b0010010100100111101000000110110110101010100111011010011001001010; end
            14'd14065 : begin out <= 64'b0010000010011101101010001110110000011001110111111010100101011010; end
            14'd14066 : begin out <= 64'b1010101101001010101010011110010100101011110010001010100100010111; end
            14'd14067 : begin out <= 64'b0010101010111111001010010011110110101000010011110010100101010011; end
            14'd14068 : begin out <= 64'b1010011011001011101010001000000100100110110010100010101001111011; end
            14'd14069 : begin out <= 64'b0010100101101101101001000010111100101001111100000010101010010111; end
            14'd14070 : begin out <= 64'b1010100001111101101001010100111100101001011110011010011110110011; end
            14'd14071 : begin out <= 64'b1010011001100111100100000001000110101001001100011010010001101100; end
            14'd14072 : begin out <= 64'b1001110000011111001010011111001100100100010100111010101110101000; end
            14'd14073 : begin out <= 64'b0010011100011001101000101011111110101011011100000010010000110100; end
            14'd14074 : begin out <= 64'b1010011010111101000101010110111000100001111110001010100111100001; end
            14'd14075 : begin out <= 64'b1010011011111100101001001000110010100011010100100010101110110101; end
            14'd14076 : begin out <= 64'b0001101100001101101010111111100010101000111101101010100100011111; end
            14'd14077 : begin out <= 64'b1010010100111000101001111001101100101011011010001010010010110111; end
            14'd14078 : begin out <= 64'b1001111111101010001010100011110010101000110000100010011110011101; end
            14'd14079 : begin out <= 64'b0010100110110011001010011101110000011000001111101010100011100000; end
            14'd14080 : begin out <= 64'b0010001000101000001010000001001000101010001000011010101011100001; end
            14'd14081 : begin out <= 64'b0010011010001011101000110011001110100101000100001010001111100010; end
            14'd14082 : begin out <= 64'b0001101010110110101010100110110100101011100100101010010001101011; end
            14'd14083 : begin out <= 64'b1010100010001111101000100001110100100100111011111010100110010011; end
            14'd14084 : begin out <= 64'b0010100001110011001000100101100000101001101110011010010001100010; end
            14'd14085 : begin out <= 64'b0010011011011011101010100101010110101000100000001010010001011101; end
            14'd14086 : begin out <= 64'b1010100101111110101000110001110000011000110111010001001110111011; end
            14'd14087 : begin out <= 64'b1010010111100010001010010011000000100001101110110010101011000111; end
            14'd14088 : begin out <= 64'b1010100100011000000101010100010000101011001101110010100000000011; end
            14'd14089 : begin out <= 64'b1010100101011011101010001111101100010100011001000010101100100110; end
            14'd14090 : begin out <= 64'b0010101010000111001001001001011010101000101010001010100111110011; end
            14'd14091 : begin out <= 64'b0010100100111100101001100111011110101001101000100010101101110100; end
            14'd14092 : begin out <= 64'b1010100111111000101010110101110010101010111100011010001100011100; end
            14'd14093 : begin out <= 64'b1010101010011011001010010000010100100011001101001010100001101110; end
            14'd14094 : begin out <= 64'b0010100110111010100111100000110100101001001011001010100100111101; end
            14'd14095 : begin out <= 64'b0010010000100001101001000001010000100101111010110010100001111100; end
            14'd14096 : begin out <= 64'b1001111101010110001010001001000100100010100111001010100011110000; end
            14'd14097 : begin out <= 64'b1010101011100011001001110010001110101001110010011001111101100100; end
            14'd14098 : begin out <= 64'b0010100010111111101010101101111010101000010111010001111010101110; end
            14'd14099 : begin out <= 64'b0010100111101000101010100110011100101000110100011010101111111111; end
            14'd14100 : begin out <= 64'b1010101110111111101000010000110110101000100010001010101000010010; end
            14'd14101 : begin out <= 64'b1001010100110111101010110001110100011010110001000010101101011101; end
            14'd14102 : begin out <= 64'b0010101001011100001000000001100100101011111111111010101110111001; end
            14'd14103 : begin out <= 64'b1010001110011111001001111010110000100111001101111010101110000100; end
            14'd14104 : begin out <= 64'b1010100101100001001010100001001100101000011100000010100111001010; end
            14'd14105 : begin out <= 64'b1010000111000111001001011001001000011100111011010010100110000001; end
            14'd14106 : begin out <= 64'b0010110000001111001010101000010010101011010100100010010101100010; end
            14'd14107 : begin out <= 64'b1010010010111100101001100010001100011011101101100010011010001001; end
            14'd14108 : begin out <= 64'b0010100000100110001010101001100100101011010101010010011010111110; end
            14'd14109 : begin out <= 64'b0010011011101010100110111000100000101011000110011010101101110110; end
            14'd14110 : begin out <= 64'b0010101110111110001010100110010010100101001111111010101010011111; end
            14'd14111 : begin out <= 64'b0010101010100111001000110001001010101000100111100010100101000111; end
            14'd14112 : begin out <= 64'b1001111110101101101001100111101110101000010001100010101010110011; end
            14'd14113 : begin out <= 64'b1010100010010011101000110000111110101011011000011010001000101011; end
            14'd14114 : begin out <= 64'b1010011101101110001010011100111000011010011101011001110110111000; end
            14'd14115 : begin out <= 64'b0010000101101110001001100111111000101010001000110001000001110010; end
            14'd14116 : begin out <= 64'b1010000000001100101010011011000110100110000011001010100100010100; end
            14'd14117 : begin out <= 64'b1010101001111010001010010011011100101001100011101010001110000100; end
            14'd14118 : begin out <= 64'b0010101110010111101010100101010010011101110010000010101110001001; end
            14'd14119 : begin out <= 64'b0010011111111001101010110010110100101011000101100010101110110001; end
            14'd14120 : begin out <= 64'b1010100100110011001001000110111010101000001011000010101011111101; end
            14'd14121 : begin out <= 64'b0010101001111110101010101001101100101000111101001010001000001100; end
            14'd14122 : begin out <= 64'b1010001111011101101001111101100110100101000011101010100110101100; end
            14'd14123 : begin out <= 64'b0010010101001101001010110111110010101011100011001010101101001010; end
            14'd14124 : begin out <= 64'b0010101011110101100110010101100010101000010000010010000101101010; end
            14'd14125 : begin out <= 64'b0010101101101001100101001101110100101011111011100010100101001110; end
            14'd14126 : begin out <= 64'b0010101011111000001000101100111010101010011100111010100111101011; end
            14'd14127 : begin out <= 64'b0010100101111001001010011100000110101010100110001010100110111101; end
            14'd14128 : begin out <= 64'b0010100101100001000111100010000100100110110011001010001101111010; end
            14'd14129 : begin out <= 64'b1010011110000110100110101011000010101000111110111001110100011100; end
            14'd14130 : begin out <= 64'b1010101111011101101000110000011110101011011101111010011100010001; end
            14'd14131 : begin out <= 64'b1010110000101101101010001101000010100010011110101010100001010111; end
            14'd14132 : begin out <= 64'b0010100001001011101001000111101100100101110011000010100010011000; end
            14'd14133 : begin out <= 64'b1010001000110000101000101000100000101001101101010010100000100111; end
            14'd14134 : begin out <= 64'b1010011101110111001010000101101010100001010111010010010111101000; end
            14'd14135 : begin out <= 64'b1001110000001101101001111011110100101000000010101010100000111111; end
            14'd14136 : begin out <= 64'b1010100001000100101001010100111010100110101101111001110100000011; end
            14'd14137 : begin out <= 64'b1010100010110110101000000001100110100100101011111010100110110001; end
            14'd14138 : begin out <= 64'b1010101000010011001010011011100010101001010110010010101100000001; end
            14'd14139 : begin out <= 64'b1010000001111010101001111111010110100000100010001010010010001001; end
            14'd14140 : begin out <= 64'b1010001101100110101001100110101010101000111101010010000010010111; end
            14'd14141 : begin out <= 64'b1001111000111001101010110101010000101000101000001001101110100011; end
            14'd14142 : begin out <= 64'b0010100010001000001010011000100010101000100010000010011110101110; end
            14'd14143 : begin out <= 64'b0010000111111101001011000000001100100101111011011010011110111010; end
            14'd14144 : begin out <= 64'b1010011100111100101010001110000110101010101101010010101101011110; end
            14'd14145 : begin out <= 64'b1010010010000000101010000110011010101011010011111010100001110100; end
            14'd14146 : begin out <= 64'b1010011010110101001010101000100110100011110101101010000001011000; end
            14'd14147 : begin out <= 64'b0010001111111101001010110110111010101011100110100010100101000000; end
            14'd14148 : begin out <= 64'b1010101011000001001001010101001010100111001011000010101101101000; end
            14'd14149 : begin out <= 64'b1010011001001110001010111101001010101001000001000010100010101000; end
            14'd14150 : begin out <= 64'b1010101000101101001000110111100010100001011100100010011101101000; end
            14'd14151 : begin out <= 64'b1001101100111110001001011011011000101011010101010010101101101001; end
            14'd14152 : begin out <= 64'b1010010100111100001001111010110000100100001111110010100001010110; end
            14'd14153 : begin out <= 64'b1010101111110010000111001110111110101011001101010010001010111110; end
            14'd14154 : begin out <= 64'b0010100010010000001010001111000100100110100011011010101010100010; end
            14'd14155 : begin out <= 64'b1010011001111111001001010100011000101011011010000010101001000101; end
            14'd14156 : begin out <= 64'b1010010001101010100111110101000110101000001001111001110110011110; end
            14'd14157 : begin out <= 64'b1010011011111100101010101000010000100001110100001010101100110000; end
            14'd14158 : begin out <= 64'b1010101001101100100111101111100100101001011100101010100110010101; end
            14'd14159 : begin out <= 64'b1001100110001001001001101100110100100111000001100010101101110010; end
            14'd14160 : begin out <= 64'b0010101000010100001000000100011100101011111100101010100100010111; end
            14'd14161 : begin out <= 64'b0010101001101100100101001000101100101010000010111010100110000111; end
            14'd14162 : begin out <= 64'b0010011010110001001001111101111110100000011010111010101010010011; end
            14'd14163 : begin out <= 64'b0010101011010011001010100001000100011110000010111010010100010110; end
            14'd14164 : begin out <= 64'b1010101111011101000111110011011110011110101111010001111010100011; end
            14'd14165 : begin out <= 64'b1010101011000110001010010000001110101000110010011010000001111000; end
            14'd14166 : begin out <= 64'b1010100101000111001001100110000010101011010000101010101001010010; end
            14'd14167 : begin out <= 64'b1010010100001110001000110100111110101010110011110010011110110011; end
            14'd14168 : begin out <= 64'b0001101001000000101010011101110100100110001111110001100111010001; end
            14'd14169 : begin out <= 64'b1001110010011111101010011110111110001001101111100010000001101010; end
            14'd14170 : begin out <= 64'b1010011110111001001010110000110100011101100010111001101111110000; end
            14'd14171 : begin out <= 64'b0010100110101101001010001000010000101010000001000010101100010010; end
            14'd14172 : begin out <= 64'b1010100001111011001010000101110000100110101100111010100011110011; end
            14'd14173 : begin out <= 64'b1010101101100111101010111000110010101000111010110010101111110000; end
            14'd14174 : begin out <= 64'b0010101110011100101010001000100110100101110100101010100000001000; end
            14'd14175 : begin out <= 64'b0010000001000110001010111000110010100111010100101010101001100110; end
            14'd14176 : begin out <= 64'b0010100010101010101001000111101000101010001011111010100010101010; end
            14'd14177 : begin out <= 64'b0001011010010110101010010100100000101000100111001010011001101101; end
            14'd14178 : begin out <= 64'b0010011101001100101010100101001000101000100101001010100000111010; end
            14'd14179 : begin out <= 64'b1010001100110111101001110010011110011111001011000010101110100001; end
            14'd14180 : begin out <= 64'b0010000010011111001000110111001010100100010011001010101111100000; end
            14'd14181 : begin out <= 64'b0010100110011001001010011001010000101010001111110010101100100110; end
            14'd14182 : begin out <= 64'b0010101010010111001010010110110010100111101000010010101101111011; end
            14'd14183 : begin out <= 64'b1001010101111010001010110101010100101010101001011001110101110001; end
            14'd14184 : begin out <= 64'b0010100110111010101010110100010010101001000111010010101111110010; end
            14'd14185 : begin out <= 64'b0010001110101010100110011011110010100001111001100010100001011000; end
            14'd14186 : begin out <= 64'b0010101001111010001000110011011010100110101011100010010111001100; end
            14'd14187 : begin out <= 64'b0010010011101000001001110011001010100111000010001010100000010010; end
            14'd14188 : begin out <= 64'b0010100110111111001001100100011000101000100111000010001111110100; end
            14'd14189 : begin out <= 64'b1010101111001100001010000111000100011110101001011010011110011111; end
            14'd14190 : begin out <= 64'b0001110100001001000111010000001110101011110111111010000010011011; end
            14'd14191 : begin out <= 64'b1010100110111101000111100100100110100011000011001001111111110100; end
            14'd14192 : begin out <= 64'b1010011100010111101001111000111000101010101111110010011000100011; end
            14'd14193 : begin out <= 64'b0010011100001110001001101100000100010010010101011010101010110010; end
            14'd14194 : begin out <= 64'b1010101000011100101001001110110110101011011111101001110100010011; end
            14'd14195 : begin out <= 64'b0010101011111011100100101110110010011110110100000010000110000011; end
            14'd14196 : begin out <= 64'b1001110111101001101001000001000110101000101100001010100110011111; end
            14'd14197 : begin out <= 64'b1010100101011010001010100101001010101001000010001010100111110101; end
            14'd14198 : begin out <= 64'b0010010101011011001000000111101000100110011110100010011000001000; end
            14'd14199 : begin out <= 64'b1010100000110100100011111101110010100100110100001010101111111101; end
            14'd14200 : begin out <= 64'b1010010000100000101000010111001010100101110000011010101000001001; end
            14'd14201 : begin out <= 64'b0010011110001010001010010010101110101010100000111001111010100000; end
            14'd14202 : begin out <= 64'b1010100010010111000101001001101010100100010110111010100111000001; end
            14'd14203 : begin out <= 64'b1010011100111001001001001011111000101001000101001010101011011001; end
            14'd14204 : begin out <= 64'b1001010010110110101000000000010100101001100001000010101010100011; end
            14'd14205 : begin out <= 64'b1010000111111001101010111100110010100011100111100010101100101100; end
            14'd14206 : begin out <= 64'b0010101000010000001010100100111100101010101100100010011001110100; end
            14'd14207 : begin out <= 64'b0010100110010110001010101000001010101001101101101010100111011010; end
            14'd14208 : begin out <= 64'b1010100110010011101001010111101010101001011101000010011101111001; end
            14'd14209 : begin out <= 64'b1010011010001011101001010110111010100010110110001010100100001110; end
            14'd14210 : begin out <= 64'b1010100111001111101001101010101100101010000111000010011101111110; end
            14'd14211 : begin out <= 64'b1010010100001011001001011110010000101011101011101010101011111110; end
            14'd14212 : begin out <= 64'b0010100001011101001010110001001010101010010111011010011101111010; end
            14'd14213 : begin out <= 64'b1010010111100110001010101010100100101011011110100010011001110111; end
            14'd14214 : begin out <= 64'b0010110000010100101001111101000110100110101010011010101011110111; end
            14'd14215 : begin out <= 64'b0010100010101001001000101010011010101011000100110010100110010100; end
            14'd14216 : begin out <= 64'b1010101110001011001001011101011100101010111001100001110111011010; end
            14'd14217 : begin out <= 64'b1010001101110111101001110110001010100100100110011010100011101100; end
            14'd14218 : begin out <= 64'b1010100001011110100110101100000000101010101001110001110000001000; end
            14'd14219 : begin out <= 64'b1010101010100010001010010000111000101010001100011001011010010101; end
            14'd14220 : begin out <= 64'b0010100110001010000111110101100100100100101011011010010011110010; end
            14'd14221 : begin out <= 64'b1010011010100100101010011011010000100100110000010010101001111011; end
            14'd14222 : begin out <= 64'b0010100101000111101001000110000010101010100100011010010110011110; end
            14'd14223 : begin out <= 64'b1010101100111010101001110110100100011001011000101010100100011100; end
            14'd14224 : begin out <= 64'b1010101001110000101001011111001100100100011011101010100111000100; end
            14'd14225 : begin out <= 64'b1001101010100100001010111100100100101001110101010010011000111001; end
            14'd14226 : begin out <= 64'b0010011001111101101001011101101100100110110010000010001100100111; end
            14'd14227 : begin out <= 64'b0010010010011100001010010011110010100111111110101010100010000001; end
            14'd14228 : begin out <= 64'b1010100000000101001010000111111010101011011100011010010101001010; end
            14'd14229 : begin out <= 64'b1010011110100000001001010111100100101000010011110010101100000001; end
            14'd14230 : begin out <= 64'b1010100101011100001010110101010010101000111101111010001111101101; end
            14'd14231 : begin out <= 64'b0010101011001101001010110111110010011001010010100010100100001101; end
            14'd14232 : begin out <= 64'b0001110010100111101010110001000100101011111111001010010101001000; end
            14'd14233 : begin out <= 64'b1010011000011011001000100110001000100110100000111010011001100110; end
            14'd14234 : begin out <= 64'b1010000110111110101010010110101000100000111000111010100101111101; end
            14'd14235 : begin out <= 64'b0010100000111111001010001011001010100111100001101001111001001001; end
            14'd14236 : begin out <= 64'b1010011000101001101010110101001100100011000100101010101010110011; end
            14'd14237 : begin out <= 64'b0010100101010111001001110010101110101010000111111010100010010010; end
            14'd14238 : begin out <= 64'b0010010110101110001010100000110100100110011111011010101000110011; end
            14'd14239 : begin out <= 64'b0010011010101010101001000001000000101010100000000010100111010010; end
            14'd14240 : begin out <= 64'b1010001110100010000110001001010010101001101100110010011000001111; end
            14'd14241 : begin out <= 64'b0010001011001100001000100111101010101010110000100010101111000101; end
            14'd14242 : begin out <= 64'b0010010110010011001001001110100110101000111001000010011011011011; end
            14'd14243 : begin out <= 64'b0010010111110110001011000000011000101000000100101000111110011010; end
            14'd14244 : begin out <= 64'b0010100000011100101001001010100110100111011100011010100101111110; end
            14'd14245 : begin out <= 64'b0010011010101111001000101001111010100011100010100010001011101101; end
            14'd14246 : begin out <= 64'b0001100000001110101001000111101110010011001110000010011001011011; end
            14'd14247 : begin out <= 64'b1010000000100000100111101000111000100011101011101010101110101111; end
            14'd14248 : begin out <= 64'b1010011001101011101001010101010110101010010010000010101011010011; end
            14'd14249 : begin out <= 64'b0001000110101111000111101111010110011110001101110010011011000111; end
            14'd14250 : begin out <= 64'b0010101001010011101001011101000000101011001100110010101000011000; end
            14'd14251 : begin out <= 64'b1010011101000011101001101010100100100110001010010001110101011111; end
            14'd14252 : begin out <= 64'b1010001001100011001001101000011010101000100001001010101001100000; end
            14'd14253 : begin out <= 64'b1010101101010101001010010100010000101010100100101010100001110110; end
            14'd14254 : begin out <= 64'b0010101000010011101001110101111100101010011101100001100110101001; end
            14'd14255 : begin out <= 64'b0010100011000000101001101001001000100110010010101001000010100100; end
            14'd14256 : begin out <= 64'b1010011100110101101010011110011110100110101001110010101100000101; end
            14'd14257 : begin out <= 64'b1010100010001011101010001101100010100010011110111010101011100111; end
            14'd14258 : begin out <= 64'b1010011001011001101000111010001100100100101000110010101110100011; end
            14'd14259 : begin out <= 64'b0010000101101111001001111010011010011011001100100001010101010011; end
            14'd14260 : begin out <= 64'b1010010111100110101010101111011000100100100010000010100010101111; end
            14'd14261 : begin out <= 64'b0010000100001000100111101000011100100101001010010010000101010010; end
            14'd14262 : begin out <= 64'b0001110101000000101001000111011110100100110111000010101011011001; end
            14'd14263 : begin out <= 64'b1010000111000001001001000000011010101010000011111010101101010001; end
            14'd14264 : begin out <= 64'b0010101001110000101010101000000000101001001101000001100111010001; end
            14'd14265 : begin out <= 64'b0001111001101010000110011111111000101001100101000010001011101011; end
            14'd14266 : begin out <= 64'b1010010100000110001001101001100110101010100011100010010001111001; end
            14'd14267 : begin out <= 64'b1010001010100011101010101001010110100100101100001010101100011101; end
            14'd14268 : begin out <= 64'b1010100101110001101010011010000100100101010101110010101000010011; end
            14'd14269 : begin out <= 64'b1010010000010111001001010110100000011111011110010010100101000001; end
            14'd14270 : begin out <= 64'b0010011100100101101010110111110100101010010100100010101111111011; end
            14'd14271 : begin out <= 64'b1010001110000100101010001110011110101001100011000001111001101101; end
            14'd14272 : begin out <= 64'b1010100101001000101001111101101100011101010110001010011111100111; end
            14'd14273 : begin out <= 64'b0001110000111110101010000110101110100001000110000010100000101101; end
            14'd14274 : begin out <= 64'b1010101000010101101010111100000000010111000011011010100110001100; end
            14'd14275 : begin out <= 64'b0010100101110110101000101001000000101001000110010010100000001100; end
            14'd14276 : begin out <= 64'b0010100010100000001010001111010100011110010011011010101011011111; end
            14'd14277 : begin out <= 64'b0010100000111100001010100101010100101000101010011010101110101001; end
            14'd14278 : begin out <= 64'b0001110101111110101001001101001010100111000100101010101011000111; end
            14'd14279 : begin out <= 64'b0001111110001010001010000010101100100010100010011010011100100100; end
            14'd14280 : begin out <= 64'b0010001000110010001010101010000100100000010111100000111110000100; end
            14'd14281 : begin out <= 64'b1010100111110101001010111011001100100101110100001010101111000101; end
            14'd14282 : begin out <= 64'b1010010011001010101000110000110000011101111011100010010001001010; end
            14'd14283 : begin out <= 64'b1010101111000101001010001000110110101011110010011001111001101100; end
            14'd14284 : begin out <= 64'b0010010011001101001010000100000000101000001011011010101110011100; end
            14'd14285 : begin out <= 64'b1010000110001011000111110000111110011101100110100001010100011000; end
            14'd14286 : begin out <= 64'b1010100111110110100111010100001000101000010010101010100101001100; end
            14'd14287 : begin out <= 64'b1010010001111110101000010101000110101011110011011010101011111101; end
            14'd14288 : begin out <= 64'b1010101110001010001010101111101110101001110111011010011101100001; end
            14'd14289 : begin out <= 64'b1010101100110100101001100111101100100100011010101010101000111001; end
            14'd14290 : begin out <= 64'b0010011000101010101010111011110100101010010001000010101111110000; end
            14'd14291 : begin out <= 64'b0010100100100111101010100110101010101001101011001010101000110001; end
            14'd14292 : begin out <= 64'b1010100010000011001010001011010100101011010011010010100010101010; end
            14'd14293 : begin out <= 64'b0010010011100000001010001100000010000110101011011010101100110100; end
            14'd14294 : begin out <= 64'b1010100101000000101010110010010100101001011001100010010011000000; end
            14'd14295 : begin out <= 64'b1010101111101010000111100111101100101001001000111010101000011111; end
            14'd14296 : begin out <= 64'b0010100011110001101001101011101000100101101100001010010010011011; end
            14'd14297 : begin out <= 64'b0001101110001000001010111000110010101010110100100010100011110110; end
            14'd14298 : begin out <= 64'b1010010001101100100110011010110110100100010101100001010011000100; end
            14'd14299 : begin out <= 64'b1001110111001111101001101000100000101010110001011010100100101111; end
            14'd14300 : begin out <= 64'b1010100000101101101010110110000100100110010100000001011111111010; end
            14'd14301 : begin out <= 64'b1010010011110111001010011110011110100111010000110010101110001101; end
            14'd14302 : begin out <= 64'b1010101011111000101001100100111010100010101010110010011011000001; end
            14'd14303 : begin out <= 64'b0010101010101101001001111100110000100101001000111010011101001011; end
            14'd14304 : begin out <= 64'b1010100101101101001000000000000110101011011100000010100011111001; end
            14'd14305 : begin out <= 64'b0010010100010001001001110001011000101010010000111010000001111101; end
            14'd14306 : begin out <= 64'b1010010011100111101010000101001110011011010100101010101110010100; end
            14'd14307 : begin out <= 64'b0010001001111111001010100011100100101011100111011010100010111011; end
            14'd14308 : begin out <= 64'b0001111110000001101010101000001110100100100110010010101000111100; end
            14'd14309 : begin out <= 64'b1010010000010100101010100110000110101001100001100010101101010110; end
            14'd14310 : begin out <= 64'b1010010111100000101010111101110110101010001100010010101000011001; end
            14'd14311 : begin out <= 64'b1001100100101101001010000110100110101000111101100010011000000100; end
            14'd14312 : begin out <= 64'b0010101111111000101000111111111100100101001101000010010110100011; end
            14'd14313 : begin out <= 64'b0010101000100010001010101100011100101000011001100010100010100110; end
            14'd14314 : begin out <= 64'b1001111000001101001010011000111100100111010111101010000001100101; end
            14'd14315 : begin out <= 64'b1010101111011111001010001011111010101011010010010001101011101110; end
            14'd14316 : begin out <= 64'b0010101000001100001001100011000000101010010011110010001101100001; end
            14'd14317 : begin out <= 64'b1010010001000110001000101011110110100100000001000010100010011000; end
            14'd14318 : begin out <= 64'b1010001001110011001001100100110110101011011010001010101111100101; end
            14'd14319 : begin out <= 64'b0010101010100011001010011101001010100111101000001010010110101111; end
            14'd14320 : begin out <= 64'b1010001011101101000111101100110000100100011101100010101010010110; end
            14'd14321 : begin out <= 64'b1010100111001110001010101010001100101011101111000010100110110001; end
            14'd14322 : begin out <= 64'b1010100101110101000110001000110000101011010101011010100001111000; end
            14'd14323 : begin out <= 64'b0010100111011101000101010101100000100111000000101010100000011110; end
            14'd14324 : begin out <= 64'b1010010010001011001010000011001010100001110010000010011100100101; end
            14'd14325 : begin out <= 64'b0010011010011010001001110011101110101011000111001010010011110011; end
            14'd14326 : begin out <= 64'b0010100001101100001000011010000100101000111010000010011111100001; end
            14'd14327 : begin out <= 64'b0010000111001010000010010111001000101001100000000001110001101111; end
            14'd14328 : begin out <= 64'b1001110001101100001010110111110100011011110011101010011101001111; end
            14'd14329 : begin out <= 64'b0010101100110011101001011100000010011000110000110010100010001100; end
            14'd14330 : begin out <= 64'b0001110101111000001010111011000000100010100100001001100110100101; end
            14'd14331 : begin out <= 64'b1010100100010001100100001100101100100100100110100010100110001111; end
            14'd14332 : begin out <= 64'b1001001110100100101001110101001000100101010010000010100101101001; end
            14'd14333 : begin out <= 64'b1010011000011111101001011001000110101000101011111001101001000101; end
            14'd14334 : begin out <= 64'b0010101010100111101010100101000010100111010100111010100001101010; end
            14'd14335 : begin out <= 64'b1010100110001000101000101100101000100111010010011001001110101000; end
            14'd14336 : begin out <= 64'b0010000001111111101001100111011100011110101001101010101100010100; end
            14'd14337 : begin out <= 64'b0010011100100001101010001100011000100111011001010010100111000111; end
            14'd14338 : begin out <= 64'b1010101000010101100110111111110000101010011101001010101110110100; end
            14'd14339 : begin out <= 64'b1010101010100001101010111111011010101011000000100010011110101000; end
            14'd14340 : begin out <= 64'b1001010011001010101010011100101010100001101111011010010001000011; end
            14'd14341 : begin out <= 64'b1010101100100100101010100101011000101010001010010010100000110011; end
            14'd14342 : begin out <= 64'b0010001011110101101001100111101000100000011111011010101110111000; end
            14'd14343 : begin out <= 64'b0010101010110011001001100000000000011010101010100010100111000100; end
            14'd14344 : begin out <= 64'b0010000110110101001000101001101000101001011100010010101101011101; end
            14'd14345 : begin out <= 64'b0010100100011101100101011101011100011110101011010010101001100101; end
            14'd14346 : begin out <= 64'b1001111000010110001000010010100010101001100001100010100010000111; end
            14'd14347 : begin out <= 64'b1010101100000001001001001110011100101000101101111010010000100111; end
            14'd14348 : begin out <= 64'b0010011100001011101010100001011010101001000111110010101111011100; end
            14'd14349 : begin out <= 64'b0010101001001010001010101101001000011100011000001010101010001011; end
            14'd14350 : begin out <= 64'b0001111011011011101010110010110110100100110001111010010110011001; end
            14'd14351 : begin out <= 64'b0010101110001101001001000000000110101010110001111001000110011000; end
            14'd14352 : begin out <= 64'b1010000001001010001010100010110100101001001001110001011101111101; end
            14'd14353 : begin out <= 64'b0001011101011010001010001101111000101001000101110010100110111011; end
            14'd14354 : begin out <= 64'b1010000101100010000111010011100100101001010101011010101110110000; end
            14'd14355 : begin out <= 64'b0010100010010011101001011100000010011111001111011001111011000100; end
            14'd14356 : begin out <= 64'b0010011111001111101010011110100100100101101100111010100011010010; end
            14'd14357 : begin out <= 64'b1010010000110101001010100010011110101010100101111010011101010100; end
            14'd14358 : begin out <= 64'b0010100011111001001001110100011010101010111100111010011100000111; end
            14'd14359 : begin out <= 64'b1010100011100101001010101001010010101000111101010010010010101110; end
            14'd14360 : begin out <= 64'b1010101100100010101010000010100010101011111011010010101111001000; end
            14'd14361 : begin out <= 64'b0010100110011111100101111001110110101000000011100010101001010000; end
            14'd14362 : begin out <= 64'b1010001111001011001010111100011110101001001110100010011110000001; end
            14'd14363 : begin out <= 64'b1010010100011110101001001000000000100101000101011010101000100000; end
            14'd14364 : begin out <= 64'b0010100100111000101010110111100100101011111001001010011001011111; end
            14'd14365 : begin out <= 64'b1001111001100101001001010110100000011111111011111010101110111100; end
            14'd14366 : begin out <= 64'b1001110011100001100111010001101100100000001111001010101100010010; end
            14'd14367 : begin out <= 64'b1010101001111011101001101001000000101010101111111010100111000100; end
            14'd14368 : begin out <= 64'b1001111011101001001010100011010000100111001000101010011101110011; end
            14'd14369 : begin out <= 64'b0001110000100001001010100010100110100110010100001010100000101001; end
            14'd14370 : begin out <= 64'b1010100000110001101010000011001010100100010001110010100000111111; end
            14'd14371 : begin out <= 64'b0010101111100101001010011100110010101000101101111010100110001101; end
            14'd14372 : begin out <= 64'b0010101101011010001010000111010100101001011100100010101010010110; end
            14'd14373 : begin out <= 64'b0010100011001010000111111010001100100110001111001010100111000111; end
            14'd14374 : begin out <= 64'b1010010111010110100110101011110010100110110000011001101100010000; end
            14'd14375 : begin out <= 64'b0010100100101100101001101001011110101000111011110010101100110011; end
            14'd14376 : begin out <= 64'b0010010001110100101001011101010000101010111100101010101001001010; end
            14'd14377 : begin out <= 64'b0010011011100111001010010001000010011110111000010010101101000001; end
            14'd14378 : begin out <= 64'b1010010110110001101001011111010010011110101011101010100111111110; end
            14'd14379 : begin out <= 64'b1010100100111100101000010110111000101000000001110010100101111111; end
            14'd14380 : begin out <= 64'b1010010000111001001001110100111010101011001001111010100110001010; end
            14'd14381 : begin out <= 64'b1010100101001010000111110110011100100111110001010010001100101000; end
            14'd14382 : begin out <= 64'b1010010100110001001001100101100010011110011101010010101110100011; end
            14'd14383 : begin out <= 64'b1010100100110010001010000100111000101010101110011010001111010111; end
            14'd14384 : begin out <= 64'b0010001101110111101001011000101010101011010011000010100011001011; end
            14'd14385 : begin out <= 64'b1010100100011010100110010010001100101011111110101010010100110011; end
            14'd14386 : begin out <= 64'b0010001100001011100101000010010000000000110011100001100011010011; end
            14'd14387 : begin out <= 64'b1010100111111011001001011101011110100100011100110010010000001101; end
            14'd14388 : begin out <= 64'b0010001000111101001010001011111000011000010001101010000101100000; end
            14'd14389 : begin out <= 64'b0010010100011110101010011111000010101011011100100010000100011011; end
            14'd14390 : begin out <= 64'b0010100011100111001001011001000010101001110111010010101011001001; end
            14'd14391 : begin out <= 64'b1010010101010011101010010000101100100101111111101010101000101010; end
            14'd14392 : begin out <= 64'b0010011001111010101001100000110100100001111101000001100100100011; end
            14'd14393 : begin out <= 64'b1010100101000110001000000011111110000101000000001001111011100100; end
            14'd14394 : begin out <= 64'b1010011000110111100110111110001110101001011110101010011000111000; end
            14'd14395 : begin out <= 64'b0010100011101011101010101110001010100101110111110010101110010010; end
            14'd14396 : begin out <= 64'b1010110000011000101001001100010110010010011001100001101011110110; end
            14'd14397 : begin out <= 64'b0010101101000110101010010101000100011100001010000010100011101100; end
            14'd14398 : begin out <= 64'b0010011111101011001000000001111010011101001011101010101101011000; end
            14'd14399 : begin out <= 64'b1001110111110100001010101001011110100110001110000010101111011101; end
            14'd14400 : begin out <= 64'b0010011001001111001000101001001100011111100101010010100000110110; end
            14'd14401 : begin out <= 64'b0010101010000110101000111110100100100100110001100010100100001110; end
            14'd14402 : begin out <= 64'b1010101101110011101010001101111010101010111011110010011110100010; end
            14'd14403 : begin out <= 64'b1001111001001100000110010111100000100011011100000010101100011101; end
            14'd14404 : begin out <= 64'b0010100000001100101010010010111010100010100010011010100110110000; end
            14'd14405 : begin out <= 64'b0001100010000100101001101011101000010110111011111010100010000110; end
            14'd14406 : begin out <= 64'b1010101110101000001000110000100100100101101011110010011010110101; end
            14'd14407 : begin out <= 64'b1010100101011010101001101010111110101001111000010010001100001111; end
            14'd14408 : begin out <= 64'b1010011101000111001010001000010110100100001001000010011100011110; end
            14'd14409 : begin out <= 64'b0010001100101001100111101000101100100001010001110010101001110011; end
            14'd14410 : begin out <= 64'b1010101010111010101001100110001110101011011000100010000111100001; end
            14'd14411 : begin out <= 64'b0010100010010111101001110000111100010101100010110010011110011111; end
            14'd14412 : begin out <= 64'b1010100010111100001010101100010100100101100101000010101010111100; end
            14'd14413 : begin out <= 64'b1001011110000111101000100000010000101010111100000010011110000000; end
            14'd14414 : begin out <= 64'b0010101010110100100101001100101110101000000010100010001111110111; end
            14'd14415 : begin out <= 64'b0010011011111000001010011001011000011111001111011010000101011110; end
            14'd14416 : begin out <= 64'b0010101000111100000111100011101000101001001100110010100110100100; end
            14'd14417 : begin out <= 64'b1010011001101001100110100010101100101000101110110010100001101101; end
            14'd14418 : begin out <= 64'b1010010110111000001001011001100010100110010100100010100100001000; end
            14'd14419 : begin out <= 64'b0010101010101011101010111101100000011100101100101010101111010000; end
            14'd14420 : begin out <= 64'b0010000100111100000111100011100100101000011010101010100110110110; end
            14'd14421 : begin out <= 64'b1010010100110011101001000101011100101010111110011010011011011011; end
            14'd14422 : begin out <= 64'b1001111000001011100111010110110010100101000110110010010101101000; end
            14'd14423 : begin out <= 64'b1010100000010110101010111110000000000111100111010010101110100010; end
            14'd14424 : begin out <= 64'b1010001110110100001010111011000010011100000110100001110010111011; end
            14'd14425 : begin out <= 64'b0010101000011100001010011001101010101011110000000010101111010001; end
            14'd14426 : begin out <= 64'b0010101100001111001010100100100100100101000110001010001100000011; end
            14'd14427 : begin out <= 64'b0010101110101011001010001001111110010000100010000010011110010001; end
            14'd14428 : begin out <= 64'b0010100110010001101010001011100110011000001111101010001110010001; end
            14'd14429 : begin out <= 64'b1010101101101100101010111101001000101010110111111010101001010010; end
            14'd14430 : begin out <= 64'b0010001111001110101010001000011100101010100110001010010001010000; end
            14'd14431 : begin out <= 64'b0010101110001100100111001000100000101000001100001010000010111010; end
            14'd14432 : begin out <= 64'b1001110101000010001001001101010110100001100011110010101000101010; end
            14'd14433 : begin out <= 64'b0010100010001001001010000110110100100010010010001010001011101000; end
            14'd14434 : begin out <= 64'b1010011000001000001010100111011110101011110001110010101001111001; end
            14'd14435 : begin out <= 64'b0010101010100100101010111100000110100111000111011010001000000010; end
            14'd14436 : begin out <= 64'b1010100100110010001010010100010000101000000111010010100001100011; end
            14'd14437 : begin out <= 64'b0010000101111000101010001000100010101010010110010010011101000101; end
            14'd14438 : begin out <= 64'b1010100011101000001001100000010000011100101000000010011110000001; end
            14'd14439 : begin out <= 64'b1010011101111010001010000010101100101011001001010010000010110010; end
            14'd14440 : begin out <= 64'b0010000001001011101010100100010000101001010000000001010111101000; end
            14'd14441 : begin out <= 64'b1010001010010011101001111111010000101010011011111010011010000001; end
            14'd14442 : begin out <= 64'b1001101101110111101001111101010000101001011011001010101000011010; end
            14'd14443 : begin out <= 64'b0010100100100000001010100110001010101001111001001010100100111100; end
            14'd14444 : begin out <= 64'b0010100110100010001010000010110000100000111000110010101100100101; end
            14'd14445 : begin out <= 64'b1010011100000001101001100000110110101011100101111010011011100111; end
            14'd14446 : begin out <= 64'b1010010111000101101010110000000000101000101111011010001000011100; end
            14'd14447 : begin out <= 64'b0010001011101111001001111010101100011100100100111010100110100010; end
            14'd14448 : begin out <= 64'b1010000011010000001010110001111100100100010000111010101001010001; end
            14'd14449 : begin out <= 64'b1010100000111100001000001000001110011000010111111010010101011011; end
            14'd14450 : begin out <= 64'b0010010111110110001010001110011110100100010110101010101011000110; end
            14'd14451 : begin out <= 64'b0010101101100111101010000101011000100110000100110010000010000111; end
            14'd14452 : begin out <= 64'b1010101000101000000111101000110000100110111001111010011101010110; end
            14'd14453 : begin out <= 64'b0010100100001110101010110000011000101001111110000010101001000101; end
            14'd14454 : begin out <= 64'b1001010010001100001001001101101100100001101000001010101101101010; end
            14'd14455 : begin out <= 64'b1010110000010100001000001110111100011101000101100010101010111100; end
            14'd14456 : begin out <= 64'b1010010010001100101000111111000000100110100010010010100010000101; end
            14'd14457 : begin out <= 64'b1010101001110110101001101011110110100110000100011010001101000111; end
            14'd14458 : begin out <= 64'b0010011010101001100111001010100100101000110100010001111111100010; end
            14'd14459 : begin out <= 64'b1010101100110110101001000101111010101001100101100010101100101100; end
            14'd14460 : begin out <= 64'b1010101101010101101010010011101010100011110000111010101010011101; end
            14'd14461 : begin out <= 64'b1010100011011001101010110011100100100111000101010010011101001010; end
            14'd14462 : begin out <= 64'b0010100011000010000110000110101010101000010001110010001111011111; end
            14'd14463 : begin out <= 64'b1010100101011100101000001111100000101001001111101010100101100101; end
            14'd14464 : begin out <= 64'b0000111000011110001000110100001010101011010110011001111010010101; end
            14'd14465 : begin out <= 64'b1010010010100001101010001011110110100001111010110010100000001011; end
            14'd14466 : begin out <= 64'b1010010111000010001000111001110010101011001110011010101001100000; end
            14'd14467 : begin out <= 64'b0010101000101010101010000110010000101001010101000001111110011111; end
            14'd14468 : begin out <= 64'b0010101110010010001010110110000010101001000101010010011100011000; end
            14'd14469 : begin out <= 64'b1010010111000001001010010110000100101011001110111010101011111111; end
            14'd14470 : begin out <= 64'b1010010011000100001010101011100110100101101011100010011110110001; end
            14'd14471 : begin out <= 64'b0010101010111100101010111111000000101000011011101010100011111001; end
            14'd14472 : begin out <= 64'b0010100000100100001001010100000100101011000101011010101111000100; end
            14'd14473 : begin out <= 64'b1010000011000011101010101001011000101011011111100010010000011111; end
            14'd14474 : begin out <= 64'b0010101101010010101010110000010100100101110110001010011110010110; end
            14'd14475 : begin out <= 64'b1010010101001110101010010011001110100100110010011010101011011010; end
            14'd14476 : begin out <= 64'b0010100001011011001010011110011100011000111100100010100011001000; end
            14'd14477 : begin out <= 64'b0001100101001100001001110100010010100001011011100010100100101010; end
            14'd14478 : begin out <= 64'b0010100100110010101001101011101110100101010000011010100011110110; end
            14'd14479 : begin out <= 64'b0010100000000000101001011001011110101010100111111010101100111111; end
            14'd14480 : begin out <= 64'b1010101101001100101010000001100010100111001101011010100110010101; end
            14'd14481 : begin out <= 64'b1010011010010011000111001111110010100110110100001010100000111000; end
            14'd14482 : begin out <= 64'b1010101011110010000101001101101000100100111011111010101010111000; end
            14'd14483 : begin out <= 64'b0001111001011000101001110000110110100111111111100010101011000001; end
            14'd14484 : begin out <= 64'b0010110000000101101010001110101100100111111100010010001111011000; end
            14'd14485 : begin out <= 64'b1010010100101011001001100000010000101010001111110010101101010011; end
            14'd14486 : begin out <= 64'b1010001001101011001010001111100100101001001001010010101110100110; end
            14'd14487 : begin out <= 64'b1010101110111100101001100011110100100100111010001010010110010010; end
            14'd14488 : begin out <= 64'b0010101010001110001010010000001100011101100011111010011011001000; end
            14'd14489 : begin out <= 64'b0010100010010110101010001001110000100101100000101010101001100100; end
            14'd14490 : begin out <= 64'b1010011000101100101010100110100000101001011110000010000011111001; end
            14'd14491 : begin out <= 64'b0010011110010000001000100010100110100000111110000010000110001100; end
            14'd14492 : begin out <= 64'b0010010001001110001001000101100010101010010001111010101000011001; end
            14'd14493 : begin out <= 64'b1010100111000010101001110100101100101010100010000010010000111011; end
            14'd14494 : begin out <= 64'b0010001011110110001010111101011010100101011000111001011000111101; end
            14'd14495 : begin out <= 64'b0010100110010111101001100010111100100111011110011010101001011101; end
            14'd14496 : begin out <= 64'b1010101001000001101001000010000100101010101101101010100010011110; end
            14'd14497 : begin out <= 64'b0010101010100001101010100010110100100011101111111010100011110000; end
            14'd14498 : begin out <= 64'b0010100111100010001001100110111100100111101001000010101100000000; end
            14'd14499 : begin out <= 64'b1001001000100011101000000110001100101011101110100010011100001010; end
            14'd14500 : begin out <= 64'b0010100110110101101001100000000010100111010010000010010000001000; end
            14'd14501 : begin out <= 64'b0001111111000100101010001001101000100111111001100010100111111111; end
            14'd14502 : begin out <= 64'b0010101100010011101010100000001110011010000011101010101100101001; end
            14'd14503 : begin out <= 64'b1010100000111111000110111010011110100100110001110010010110011100; end
            14'd14504 : begin out <= 64'b0010101110100011000111001100110100100010101001011010010101101100; end
            14'd14505 : begin out <= 64'b1010011000111001101010010110000000101001001011110010100101001000; end
            14'd14506 : begin out <= 64'b0010011101111110000111110011110010101010001010001010010101111101; end
            14'd14507 : begin out <= 64'b0001010100010100101000110000100010100101110010101001011000000101; end
            14'd14508 : begin out <= 64'b0010000000101000001001100110010100100110001010101010011110001101; end
            14'd14509 : begin out <= 64'b0000111000001110101010101101100100011000101011101010100011011001; end
            14'd14510 : begin out <= 64'b1010010000101000001010100110100000100100000100101010101010111110; end
            14'd14511 : begin out <= 64'b0010000111111111101010000010101010101000011011011010011111010010; end
            14'd14512 : begin out <= 64'b0010011011001011001010011101111000101010100110110010010010011000; end
            14'd14513 : begin out <= 64'b1010010001101111101001011101011000100001100010011010100010000000; end
            14'd14514 : begin out <= 64'b1010100101101110101001011111010010101001101101111010101110111110; end
            14'd14515 : begin out <= 64'b1001110101001111001001011000000100100001111100110010100000000011; end
            14'd14516 : begin out <= 64'b1001111010110110101001010110001000100101101011111010011010000111; end
            14'd14517 : begin out <= 64'b0001100111110101001001101011100100100001011100100010010001001001; end
            14'd14518 : begin out <= 64'b0010101000011101001010011000111000011010010000111001110001011001; end
            14'd14519 : begin out <= 64'b0010100100000011101010111010001110101000000001110010101111000010; end
            14'd14520 : begin out <= 64'b1010010000011110100110001011111000100100111010010010001010110010; end
            14'd14521 : begin out <= 64'b0001110000011000001010001001110100101010001111100010100000010110; end
            14'd14522 : begin out <= 64'b0010100010011100101010111100110000101000110000110010001010111000; end
            14'd14523 : begin out <= 64'b1010011101101001101010101011111100101000100110111010100010100010; end
            14'd14524 : begin out <= 64'b0010001101100101101010110101001100101011010011000010101111001011; end
            14'd14525 : begin out <= 64'b0010101110100000001010011100010100101000001011110010001000011101; end
            14'd14526 : begin out <= 64'b1010100011011111101001011101101110100111111001010001110011010111; end
            14'd14527 : begin out <= 64'b0010001110001000101001111101100100001100011011100010001010111001; end
            14'd14528 : begin out <= 64'b1010100000101011001001101110101110100001011100000010101010100000; end
            14'd14529 : begin out <= 64'b0001001011111001001010111010100000101010010011110010100110010110; end
            14'd14530 : begin out <= 64'b0010100000100001101010101100011100100011100101011010011100100111; end
            14'd14531 : begin out <= 64'b0010010000100101001001010010000000100111101110000010100100011010; end
            14'd14532 : begin out <= 64'b1010101010000101001010000011001010101001011101011010101111001100; end
            14'd14533 : begin out <= 64'b0010101110110011001010001010001110010101111100111010100011101000; end
            14'd14534 : begin out <= 64'b0010101100000101001000010000111110101001110111000010100010101111; end
            14'd14535 : begin out <= 64'b0010011101110110101010001001010110100111111010011010101110111110; end
            14'd14536 : begin out <= 64'b1010101100111001001010001010011000101011001111100001100001101101; end
            14'd14537 : begin out <= 64'b0001010001111011101010100000000100011101000100010010101110010001; end
            14'd14538 : begin out <= 64'b0001110100101101101000111110010010101011110110111001110110011011; end
            14'd14539 : begin out <= 64'b1000111001101011001010001001011100101000000010011010011010101001; end
            14'd14540 : begin out <= 64'b0010100000100110001010101010110010100100000100101010100111010111; end
            14'd14541 : begin out <= 64'b0001111110001001101001101010100000101010010100111001000011001100; end
            14'd14542 : begin out <= 64'b0010101011111010101010010000011100101001001010111010001000010100; end
            14'd14543 : begin out <= 64'b0010011000110110000101010111100010100010100011110010010010011111; end
            14'd14544 : begin out <= 64'b1010011110010001001010001010001110101010101011010010000011111001; end
            14'd14545 : begin out <= 64'b0010010001100010101010010100000010100000000100000010001111100101; end
            14'd14546 : begin out <= 64'b1001101110000000001010001110000010100100111111101010100000001100; end
            14'd14547 : begin out <= 64'b0010001010011010101000000011100100101001011100011010101001011011; end
            14'd14548 : begin out <= 64'b0010001111000101101001110111110110101010111101000010010011001111; end
            14'd14549 : begin out <= 64'b0010101111010001101010101011011110011110100111000010101110001001; end
            14'd14550 : begin out <= 64'b0001110010001100001000010011100100101010000010001010100101011001; end
            14'd14551 : begin out <= 64'b0010100001001000101010011111000110101001111110100010101011000101; end
            14'd14552 : begin out <= 64'b1010100110100101001010101000111110101000111101111010010001001011; end
            14'd14553 : begin out <= 64'b0010101110001000001010100101100100101010011101110010100100001110; end
            14'd14554 : begin out <= 64'b0010011101100011000111101100110010100101011000110010000000101011; end
            14'd14555 : begin out <= 64'b0010101001011000101010000000101000101001101001010010101000011001; end
            14'd14556 : begin out <= 64'b0010011101000001101010011001111110101000110011010010100000101111; end
            14'd14557 : begin out <= 64'b0010101110000101001001010011100010101000001110110010101111111000; end
            14'd14558 : begin out <= 64'b0010010011001100001010001101100110100001001001001010101111000001; end
            14'd14559 : begin out <= 64'b0010101010001101001010101001111100011100001010011001100001000000; end
            14'd14560 : begin out <= 64'b0010100001010011001010010110000110100101011110111010100000000111; end
            14'd14561 : begin out <= 64'b1010100000011001001001001000011010101010110011100010101000111010; end
            14'd14562 : begin out <= 64'b0010100010100001001010011100101110100110001111110000110000000011; end
            14'd14563 : begin out <= 64'b0001110110100110101000101011101100101001110010010010011100010100; end
            14'd14564 : begin out <= 64'b0010100110100000001001001010010010010101101101100010101010011001; end
            14'd14565 : begin out <= 64'b1010100010110111101010110100110010011101111110100010000001000010; end
            14'd14566 : begin out <= 64'b0010001111111101001010100001000000100111111111010010101111101100; end
            14'd14567 : begin out <= 64'b1010010110011110101010010110001010011110001001011010100011011100; end
            14'd14568 : begin out <= 64'b0010101001000000101001010000011010100001111001000001011010001000; end
            14'd14569 : begin out <= 64'b0010010101101101101010011110010110101000000111111001111101010110; end
            14'd14570 : begin out <= 64'b1010100000010110001010100010101010100010111100100010100000110000; end
            14'd14571 : begin out <= 64'b0010011101110000001010100110000010100000110111011010001100000110; end
            14'd14572 : begin out <= 64'b0010100001101100101000000010001000101001000100000010100101100000; end
            14'd14573 : begin out <= 64'b0010000000010011101010010010001010010101010010111010000010110000; end
            14'd14574 : begin out <= 64'b0010010010011001001010101010110110100010100111110010000001000101; end
            14'd14575 : begin out <= 64'b0010101010000001101010110100110010100001100101000010100010000100; end
            14'd14576 : begin out <= 64'b1010011000111011101000000101011110100101110111110010100110001101; end
            14'd14577 : begin out <= 64'b0010101101111101001010111111100000100000111100111001001000101110; end
            14'd14578 : begin out <= 64'b0010101010010111101001001110101110100011111110111010100000100111; end
            14'd14579 : begin out <= 64'b0010000111111001101010011110001010100101110111011001111110011110; end
            14'd14580 : begin out <= 64'b1010001010011101101010101111010110100110010011011010101111101000; end
            14'd14581 : begin out <= 64'b0010000000010111101010111011111000100101100100010010011110000101; end
            14'd14582 : begin out <= 64'b1010101101101101001001100010001100101000110111101010011110111111; end
            14'd14583 : begin out <= 64'b1010100000000000101010100011000110100100001110011010001100001101; end
            14'd14584 : begin out <= 64'b0010101101100110101010000111101000101010000111011010011100001100; end
            14'd14585 : begin out <= 64'b0010100011111110101001000011010100101000011010000010101110100100; end
            14'd14586 : begin out <= 64'b1010000101101110101000101100011010101000100101001010010110101111; end
            14'd14587 : begin out <= 64'b0010100110001111101010111011101010100011010001010001101000000011; end
            14'd14588 : begin out <= 64'b0010011101011110001000111000010100011111100001101010101111101111; end
            14'd14589 : begin out <= 64'b0010100100110110101000111101011000101010010010000010100110011011; end
            14'd14590 : begin out <= 64'b1010001101001101001010000011000000101010011010111001100100100100; end
            14'd14591 : begin out <= 64'b1010101011010110001010110111010000101000101010001010101000010000; end
            14'd14592 : begin out <= 64'b1010101101000000000111000000011000100000101010010010001010101110; end
            14'd14593 : begin out <= 64'b0010011100100101101001011101011100010000101100100010100001010101; end
            14'd14594 : begin out <= 64'b0010101110010101101010111001111010101000101000011010101100100001; end
            14'd14595 : begin out <= 64'b1010000101110010001010101111101110101000000100110010101110111001; end
            14'd14596 : begin out <= 64'b1010001101011101100110101011101000100110010111110010010010011011; end
            14'd14597 : begin out <= 64'b0001110100000100001010011001011110100000110011011010000000011001; end
            14'd14598 : begin out <= 64'b1010010111110101101000001100001110100010111101001010100111100011; end
            14'd14599 : begin out <= 64'b1010100000101101100111100001001010100010000011100010100001101011; end
            14'd14600 : begin out <= 64'b0010101111011101101001101011110110011101000010010010101111101111; end
            14'd14601 : begin out <= 64'b0010100101111111001001011010010100101100000011011010100101101110; end
            14'd14602 : begin out <= 64'b1010100011111000001010010101101010101010011100100010101110010001; end
            14'd14603 : begin out <= 64'b1010010000110011101010000100100010101000010011000010100110010111; end
            14'd14604 : begin out <= 64'b1010011001110000100111100100000000101001010011000010100111000010; end
            14'd14605 : begin out <= 64'b1010100011100111100111000100111100101011100010110010000001111110; end
            14'd14606 : begin out <= 64'b1010101000000001000110011010111100101001111111100010110001011110; end
            14'd14607 : begin out <= 64'b1010100010101000001010000101111010101011101000110010101111100100; end
            14'd14608 : begin out <= 64'b1010101011101100001010110010001100100110000101110010010001001111; end
            14'd14609 : begin out <= 64'b1010010110101101001001101110111100101010101010110010010100000011; end
            14'd14610 : begin out <= 64'b0010000001100010100011011011000000100001010000110010101110100010; end
            14'd14611 : begin out <= 64'b1010010110001110001010011110110010101000101100010010101000111011; end
            14'd14612 : begin out <= 64'b1010011110111001001010010010110110101010011100101010000001010100; end
            14'd14613 : begin out <= 64'b1010101010110100001010111110111010101010101111010001111100111111; end
            14'd14614 : begin out <= 64'b0001111010000011101010011000001100011000001010011010101100111110; end
            14'd14615 : begin out <= 64'b0010101010001110101010011001101000101001001001100010110000001111; end
            14'd14616 : begin out <= 64'b0010100111011110001000110010100110100110000010100010100011101110; end
            14'd14617 : begin out <= 64'b1010100111100111001010010000000100101001101001010010101100111111; end
            14'd14618 : begin out <= 64'b0001011110110101101001110000100100101001111010111001111010110010; end
            14'd14619 : begin out <= 64'b0010101101101001001010111101011010101001110000000010101100010010; end
            14'd14620 : begin out <= 64'b0010101000001111100111000000001010101011111010001010101011000110; end
            14'd14621 : begin out <= 64'b0010100000101000101010000011000010100000000011110010100010011100; end
            14'd14622 : begin out <= 64'b1010010000011010000111000010110110101000111111011010100101100011; end
            14'd14623 : begin out <= 64'b1010011000011000101010100010000000101001011000100010101100001111; end
            14'd14624 : begin out <= 64'b1001111011101101001010101111111100100111110111001010100011101101; end
            14'd14625 : begin out <= 64'b1001110011101000101001000000001110011101001001111010101100110110; end
            14'd14626 : begin out <= 64'b1010011001001010001010111010100010001100101000010010101001011100; end
            14'd14627 : begin out <= 64'b1010000010111001001000110111000010101001010110010010100111111100; end
            14'd14628 : begin out <= 64'b0010010011000010101010101010100100101000011111000010010101110111; end
            14'd14629 : begin out <= 64'b0010001110000000001010011001011100010111001000111010101100100010; end
            14'd14630 : begin out <= 64'b1010101110100101001001000110101000101000010101010010010001101111; end
            14'd14631 : begin out <= 64'b1010100111000111001010111111100000100011110110111001101101110100; end
            14'd14632 : begin out <= 64'b1010101111010101001001100101011000011110111111111010101010101010; end
            14'd14633 : begin out <= 64'b0010010100010010001010000001001010100111110001001010100000011000; end
            14'd14634 : begin out <= 64'b0001011110001010001001101000110010101000110001101010010001010000; end
            14'd14635 : begin out <= 64'b1010101110110101001001100100001110100111001011110010010000101100; end
            14'd14636 : begin out <= 64'b1010100000110111001010000101111100100000011011100010100011001111; end
            14'd14637 : begin out <= 64'b0010101101110000001001110011110010101011100111001010010010000001; end
            14'd14638 : begin out <= 64'b0010000110111101001000001011000100101000001111011010101001001011; end
            14'd14639 : begin out <= 64'b1010100110101001001000100101001100101000111001101010100010110110; end
            14'd14640 : begin out <= 64'b1010011001110001101001110111010010010100100111100010001100010100; end
            14'd14641 : begin out <= 64'b1010001011111110100110111111011000101001111000011010100110010110; end
            14'd14642 : begin out <= 64'b0010000011101001101001110111000010011101000100011010101111101110; end
            14'd14643 : begin out <= 64'b0001110111000010100011001100000010101100000111101010010001111000; end
            14'd14644 : begin out <= 64'b0010011111010000001000011011111000100101001011110001110101100011; end
            14'd14645 : begin out <= 64'b1010101111111101101010011010001000100010010010110010010111010001; end
            14'd14646 : begin out <= 64'b1010001010100000001001100110111010011100101010101010000010110010; end
            14'd14647 : begin out <= 64'b1010101111011101001001111110111000100101110100010010010110111001; end
            14'd14648 : begin out <= 64'b0001110000110100101010000000111000101000110110100010011010001001; end
            14'd14649 : begin out <= 64'b0010100001000110001010110000010110101001100000101010001110001000; end
            14'd14650 : begin out <= 64'b0010101111101110001001001110011010101010110011110010010011011111; end
            14'd14651 : begin out <= 64'b1010010100100001001001011111011000011001011011010010100100101001; end
            14'd14652 : begin out <= 64'b1001110110100101001000101011101110100100100111110010001001110000; end
            14'd14653 : begin out <= 64'b1010101001100011001001110101111110101011111111101000111000011100; end
            14'd14654 : begin out <= 64'b1001011111000011101010111000010110010111011010000010011110100001; end
            14'd14655 : begin out <= 64'b0010010001101000001010001101111110100010011010111010010110101001; end
            14'd14656 : begin out <= 64'b1010000100111111101010000111010100100101101010110001110011011110; end
            14'd14657 : begin out <= 64'b1010100100111110001010110011101100011111010001101010000100110111; end
            14'd14658 : begin out <= 64'b0010100010000000001001011111010100101000111100101010100100011001; end
            14'd14659 : begin out <= 64'b1010101010110101001011000000000000100001101011010001111111100100; end
            14'd14660 : begin out <= 64'b1010011010100011101000011100001010101001000110001010101010001101; end
            14'd14661 : begin out <= 64'b1010010011011100100101010000100110100101010111101010001000101010; end
            14'd14662 : begin out <= 64'b0010010010110100100111100011100110101011011011000010101001100101; end
            14'd14663 : begin out <= 64'b0010011011111001101010100100100000101000110100110001010011000000; end
            14'd14664 : begin out <= 64'b1000110100001100000111111111101000100001100000010010100111111010; end
            14'd14665 : begin out <= 64'b1010101100011100101010000100111010100111111111111010100000011010; end
            14'd14666 : begin out <= 64'b0010100001001111001010100100001010100010010011111010010001011001; end
            14'd14667 : begin out <= 64'b1010000111110011101010100001111010101010111111111010010110110101; end
            14'd14668 : begin out <= 64'b1010101010101000101010100011111000011110101011010010010101001010; end
            14'd14669 : begin out <= 64'b0010011011000101101010100001011110100111101001011010100110011000; end
            14'd14670 : begin out <= 64'b1010011010000100101010000010010110010101001110000010100111000001; end
            14'd14671 : begin out <= 64'b0010100000101101001010010110100010100110111011101010101101111111; end
            14'd14672 : begin out <= 64'b0010101111000101101001010001001000100100001000100010011011001011; end
            14'd14673 : begin out <= 64'b1010100000010010001010000001000000101000110100101010101010110011; end
            14'd14674 : begin out <= 64'b1010010110111110001001000000110110011001000000000001001011011100; end
            14'd14675 : begin out <= 64'b0010010000100001001010011101010010100011100110001010000101011110; end
            14'd14676 : begin out <= 64'b1010100010100100001001011011011000100100110100000010101001000111; end
            14'd14677 : begin out <= 64'b0010100101100110101001101000000100100100100001101010101001100011; end
            14'd14678 : begin out <= 64'b0010000110001101000100000111111000100111001100000010011101100110; end
            14'd14679 : begin out <= 64'b1010011001101101101000110111111110101001000111101010101111010110; end
            14'd14680 : begin out <= 64'b1010100110100111001001001010011100100100011101000010100001000001; end
            14'd14681 : begin out <= 64'b1000111011010111001010111000010010101010001100000010001001111000; end
            14'd14682 : begin out <= 64'b1010000000010001101010010110001100101000010100001001110110000000; end
            14'd14683 : begin out <= 64'b0010101000000110000110011101101010101011101000111000010111110000; end
            14'd14684 : begin out <= 64'b0001110101010000101001110001101110100010111110100010101100011010; end
            14'd14685 : begin out <= 64'b1010100110111101101001100001000010101001000001011010001111100010; end
            14'd14686 : begin out <= 64'b0010000000110010000111111001100110101000011101101010011101111000; end
            14'd14687 : begin out <= 64'b1001111111011010101010001001010100100101000001011010101001100000; end
            14'd14688 : begin out <= 64'b1010101110111101101010101111011100101001110101100010100001010000; end
            14'd14689 : begin out <= 64'b1010000010101001001010001010000110101000110011111010100010100001; end
            14'd14690 : begin out <= 64'b0010011010100100101010100011101010101010101011010010100000110100; end
            14'd14691 : begin out <= 64'b1010011100101000101010001001000110101001011101000010100000110000; end
            14'd14692 : begin out <= 64'b1010011000000111001001000010000010101001010010101010100001001001; end
            14'd14693 : begin out <= 64'b1010100011001111001010101100100110101011001101101010100000010110; end
            14'd14694 : begin out <= 64'b1010100111011001001010101110100110010001000111101010001111110011; end
            14'd14695 : begin out <= 64'b0001001111001110101010011010001100101010111110010001100110001010; end
            14'd14696 : begin out <= 64'b1010011101101101100111010010100110100010111101001010101001010001; end
            14'd14697 : begin out <= 64'b0010101111001110001010111111111000100001100110101010101000101001; end
            14'd14698 : begin out <= 64'b1010011011011111001010110000111110100101111110101010101100100010; end
            14'd14699 : begin out <= 64'b1010010111110001100111001111000100010011111101011010010000001101; end
            14'd14700 : begin out <= 64'b1010100110010000101010110001000000101010010010000010101001101110; end
            14'd14701 : begin out <= 64'b0010010110011001101000111101000100101000111011000010000101011000; end
            14'd14702 : begin out <= 64'b1010001001110100001001111110101110100000101111111010100110101001; end
            14'd14703 : begin out <= 64'b0010010001001100001010000010111110100111010111111010101010010010; end
            14'd14704 : begin out <= 64'b1010100100110001001010110010100000101010111010100010101011011100; end
            14'd14705 : begin out <= 64'b0010101001111001001000111111100110101011101101000010101011100011; end
            14'd14706 : begin out <= 64'b0001111110001000100100010100110110100101101101111010000100001000; end
            14'd14707 : begin out <= 64'b1010100010110101001001010010001000101000000101011010000111100100; end
            14'd14708 : begin out <= 64'b0010100010111010001001000001101110101011011110000001111011111100; end
            14'd14709 : begin out <= 64'b1010101010001000001010100100001110100101010101111010101100111010; end
            14'd14710 : begin out <= 64'b1010101100110111101000100100100100101010100100010010100001100000; end
            14'd14711 : begin out <= 64'b1001111011001011100011111101101010011111100011010010010000110100; end
            14'd14712 : begin out <= 64'b0010101000000011101010000001001100101010010011100001101000101111; end
            14'd14713 : begin out <= 64'b1001111010010111101010100011111100100101100110100010001100110001; end
            14'd14714 : begin out <= 64'b1010011000010001001010110101110010100000110010101010010001000001; end
            14'd14715 : begin out <= 64'b0010101000110000001010001010101000011011111010001010011111010010; end
            14'd14716 : begin out <= 64'b0000100001000110001010110110001100100100101011101010101010000110; end
            14'd14717 : begin out <= 64'b0001111110101111101000110000101110101011001100100010010100011010; end
            14'd14718 : begin out <= 64'b0010000110000011101010100111111000100101001011100010100111110110; end
            14'd14719 : begin out <= 64'b0010100011001010001001001100100010101011011100100010101001100010; end
            14'd14720 : begin out <= 64'b1010101010110110101010100010000010101001011101001010001110000100; end
            14'd14721 : begin out <= 64'b0010100001001011101000000111111100101100000100000010100110001100; end
            14'd14722 : begin out <= 64'b0010011111100011001001000100100010101010010101000010100101010011; end
            14'd14723 : begin out <= 64'b1010011111010011101001110110110110101010101000100010100111101011; end
            14'd14724 : begin out <= 64'b0010010000101001001001010000010100101000011000100010001010111011; end
            14'd14725 : begin out <= 64'b0010010110101010001010101000001010101011011111111010011101111001; end
            14'd14726 : begin out <= 64'b0010010011000000101010101111101110101001011100111010100011011000; end
            14'd14727 : begin out <= 64'b1010100101011100101010011111010100011111111000001010010001101110; end
            14'd14728 : begin out <= 64'b1010011110000000001001000111110000101011011001011010101000111101; end
            14'd14729 : begin out <= 64'b1010001111101101101010010001010000101011110011110010101100011110; end
            14'd14730 : begin out <= 64'b0010010100111111101001011000111010011101110110011010011100010001; end
            14'd14731 : begin out <= 64'b0010100011100111101001100110100100101011001100111010100101100000; end
            14'd14732 : begin out <= 64'b1010001100100101001010100001000000100100111011111010010001000001; end
            14'd14733 : begin out <= 64'b1010010010010110101010011101110110100000001010101010010000101111; end
            14'd14734 : begin out <= 64'b1010010111001101001010000001110010100011101011000001111000011111; end
            14'd14735 : begin out <= 64'b0010010101101100101010000000010010101011101110010010000001110100; end
            14'd14736 : begin out <= 64'b1010101101001110001010100111010110101001101000001010101111110010; end
            14'd14737 : begin out <= 64'b1010101001100101101010110011111100101000110000101010100100100100; end
            14'd14738 : begin out <= 64'b0010101111111011101010011000101010010001100101100010101000110011; end
            14'd14739 : begin out <= 64'b1010011110100001001000111001000010100111000101111010101000010100; end
            14'd14740 : begin out <= 64'b0001100000111001001001101110010100101010100101110010010000000100; end
            14'd14741 : begin out <= 64'b0001101100000001001000110101101000101010110101100010100001101011; end
            14'd14742 : begin out <= 64'b0010101010100100101001111011101110011001010101011010001100011100; end
            14'd14743 : begin out <= 64'b0010100001011111001000010111111100100111011000000010010000001001; end
            14'd14744 : begin out <= 64'b0001111000001001101010010100101000101000100110011001111001000110; end
            14'd14745 : begin out <= 64'b1010101101100110001010110001101000101000010011111010100111110011; end
            14'd14746 : begin out <= 64'b1010010001011010101000000100011110100010011000000001001111010011; end
            14'd14747 : begin out <= 64'b0010011010001111101010010110101100100100100010111010100010001111; end
            14'd14748 : begin out <= 64'b0010011010011100001010101011011110101000001110010010011000011100; end
            14'd14749 : begin out <= 64'b0010101010101010101001111000101000101001110110101010001010011101; end
            14'd14750 : begin out <= 64'b0010010111101101001010111001100000100001100100011010000101101111; end
            14'd14751 : begin out <= 64'b1010101110100101101010110100011110100100111101010001101100110010; end
            14'd14752 : begin out <= 64'b0010101010100000001000101110000010100010001011000010100011110011; end
            14'd14753 : begin out <= 64'b1001110010110100001001000000111100001000001000010010000110110111; end
            14'd14754 : begin out <= 64'b0010101110110110101010010100101100101010001001111001111101011001; end
            14'd14755 : begin out <= 64'b1010100100100110001001100000100010101010001110011010101011101000; end
            14'd14756 : begin out <= 64'b0010010100001110101010101111110110101000101111011010000010001010; end
            14'd14757 : begin out <= 64'b1010100100111101101001011011000010100101001001011001110001110011; end
            14'd14758 : begin out <= 64'b1010100101100010001010010000011100101010010011101010100010110001; end
            14'd14759 : begin out <= 64'b1010101101101101001001101010101110100101110010010010100101011100; end
            14'd14760 : begin out <= 64'b0010101011110001101001110110010010101011001111001001111101101111; end
            14'd14761 : begin out <= 64'b0010010000111010101010110101010010101011101101011010010110010111; end
            14'd14762 : begin out <= 64'b0010100000001011101001110111101010101000110101010010101101101100; end
            14'd14763 : begin out <= 64'b1010100001011110101001110111100010101000011001101010011000000100; end
            14'd14764 : begin out <= 64'b0010000111101001001010001011100010011110111110101010001001101110; end
            14'd14765 : begin out <= 64'b1010011001110010101001010000011000100101011011111010011001010101; end
            14'd14766 : begin out <= 64'b0010101011001011101001011110101000101010110001011001110011001110; end
            14'd14767 : begin out <= 64'b0010101101110010101010101111110000101001111100000000000111001010; end
            14'd14768 : begin out <= 64'b0010010100100011001010101101110010100100111001110010101010110111; end
            14'd14769 : begin out <= 64'b1010101000010101101010100001001100101000000011101010100101010101; end
            14'd14770 : begin out <= 64'b1010100110110100001011000000011000100100100110001010100010000111; end
            14'd14771 : begin out <= 64'b1010100101111010001000010001010010100101010001100010101001111101; end
            14'd14772 : begin out <= 64'b0010101100100001001010101110101110100011101110000010010110001010; end
            14'd14773 : begin out <= 64'b0010100000001011001000110111111100101011100000110010011011111111; end
            14'd14774 : begin out <= 64'b1010000100110110001010100111101000101000100010001010101100100001; end
            14'd14775 : begin out <= 64'b1010000010111000001001110110011100101001110101010010101000000001; end
            14'd14776 : begin out <= 64'b0010100100100111001010000110011110101000010011011010001010001010; end
            14'd14777 : begin out <= 64'b1010000011111010101010011101100110100111011001011010010100001111; end
            14'd14778 : begin out <= 64'b1010100011000001101000011001000000101010000101000010001011100110; end
            14'd14779 : begin out <= 64'b1010100110111010101010011001000000101000101010100010100110010010; end
            14'd14780 : begin out <= 64'b0010100111100101101010100110000110101000000000101010011000011100; end
            14'd14781 : begin out <= 64'b0001010100001100101010011010011110011111100010001010100001010110; end
            14'd14782 : begin out <= 64'b1010100010011110101001100001100110100000000000100010100011111010; end
            14'd14783 : begin out <= 64'b0010011001100110001010110110011110010111111100110010001011100000; end
            14'd14784 : begin out <= 64'b0010011010011101101001010100000100100111100001000010101000101000; end
            14'd14785 : begin out <= 64'b0001110110101000101001001111100100011011100111001001011100111100; end
            14'd14786 : begin out <= 64'b0010000001010100100111111111100010100001001000000010000001110011; end
            14'd14787 : begin out <= 64'b1010100001010000001000010111011110011110000011001001000100110101; end
            14'd14788 : begin out <= 64'b0010100001001100101000011010000000101010000011111010100101011011; end
            14'd14789 : begin out <= 64'b0010001010010010001001000000010110100100001010011010100110111010; end
            14'd14790 : begin out <= 64'b0010101011000000001010000000011000101010001000001010110000100010; end
            14'd14791 : begin out <= 64'b1010011111110000001000011010001110101000011011011010101111010101; end
            14'd14792 : begin out <= 64'b0001110000000110001001000110101010011011111001110010101000110000; end
            14'd14793 : begin out <= 64'b1010001011100110000110000111110010101010000100101010100110011001; end
            14'd14794 : begin out <= 64'b0001100011001101101010011101001000101011011101100010100101001011; end
            14'd14795 : begin out <= 64'b1010101110110001101001101011101000100101001010110010011011010110; end
            14'd14796 : begin out <= 64'b0010011111101101001011000000000000100000110010100010101000101010; end
            14'd14797 : begin out <= 64'b0010001111110111000111011001111110100011010111001010011011110000; end
            14'd14798 : begin out <= 64'b0010010110011010101001110110111010101000111011101010100110000110; end
            14'd14799 : begin out <= 64'b1010010101110100101010011101000000011111000000111010100111001110; end
            14'd14800 : begin out <= 64'b1010010001100101101010111101101100101001011101100010001010110001; end
            14'd14801 : begin out <= 64'b1010100011110010101010101010111000101010010010100010010100101010; end
            14'd14802 : begin out <= 64'b0010011001101010101000110000011100101000011100111010100100000000; end
            14'd14803 : begin out <= 64'b0010010101110111001010100000100000101000110100111010000110010000; end
            14'd14804 : begin out <= 64'b0010100100100010101010100011101100101010101010001001101000000011; end
            14'd14805 : begin out <= 64'b0010101010010000000111110001011100101010000011010010101011010110; end
            14'd14806 : begin out <= 64'b1010101101000001101001000111000000100000001101011010101011110101; end
            14'd14807 : begin out <= 64'b1010010111100010101010111101111010100000000110011010011011101110; end
            14'd14808 : begin out <= 64'b1010100100011001101010101001100100100011010111011010100001111001; end
            14'd14809 : begin out <= 64'b1010011111110011001010010000110110101001000000100010011100110010; end
            14'd14810 : begin out <= 64'b1010101001110000001010001011001000011000110001110010010111101011; end
            14'd14811 : begin out <= 64'b1010100101101001101010010000101000101010101011001010100101010011; end
            14'd14812 : begin out <= 64'b0010100100001001101000001100100010100000110110110010100000110100; end
            14'd14813 : begin out <= 64'b0010100111000101001010101011000000100011001100111010011011001010; end
            14'd14814 : begin out <= 64'b1010100101000100001001010111111000101010001101001010100000010101; end
            14'd14815 : begin out <= 64'b1010101001111111001000000110000110101011111011100010101001011001; end
            14'd14816 : begin out <= 64'b0001110110100101001010010111111010101011010100100010011111101001; end
            14'd14817 : begin out <= 64'b1010101100001011101010000111000010100001000001111010100110011100; end
            14'd14818 : begin out <= 64'b0010001010101101001010100000001010101011101011111010100010110111; end
            14'd14819 : begin out <= 64'b0010000110100100001000000010100100101010111001110010100000000000; end
            14'd14820 : begin out <= 64'b0010100110000010101010111100110010100000010000111010101100011010; end
            14'd14821 : begin out <= 64'b0010101101111111100111011101100110011001001101100010101000001110; end
            14'd14822 : begin out <= 64'b1010011101100000101001100010001000100101111011111010010010000110; end
            14'd14823 : begin out <= 64'b0010101000000110101001101011110110100011111011100010100111111110; end
            14'd14824 : begin out <= 64'b0001111011101000001000011010010100101001000101101010011000101100; end
            14'd14825 : begin out <= 64'b0010100011001100101010001000100100100011011011111010000000011100; end
            14'd14826 : begin out <= 64'b0010101011100011001000000000110000101010011010101010101100110101; end
            14'd14827 : begin out <= 64'b0010101001111010101010011010010000100111001001100010101101100010; end
            14'd14828 : begin out <= 64'b0010100001110000001011000010101100100000101011111010101000000001; end
            14'd14829 : begin out <= 64'b1010000011000010001001100101101100100101100111110001110111100101; end
            14'd14830 : begin out <= 64'b1010010100100010001010100000110110011000110101000010100001110100; end
            14'd14831 : begin out <= 64'b0010101110101101001010010011111110011100101101101010010100110011; end
            14'd14832 : begin out <= 64'b1010100100010001101001101010110100011100110001110010010000111100; end
            14'd14833 : begin out <= 64'b1001111010000000100100001100100110101000111100000010010000111010; end
            14'd14834 : begin out <= 64'b0010010000110101001010101110100010100010000010100010000010001101; end
            14'd14835 : begin out <= 64'b0001000111010100000110010110100100101011010011101010101110111101; end
            14'd14836 : begin out <= 64'b1010101110001110001000000110001010101000001010011010100100001111; end
            14'd14837 : begin out <= 64'b1010001111101010101001100011001000101010000001001010001011011011; end
            14'd14838 : begin out <= 64'b0010100010101011001010111110111000101010100001011010011101001010; end
            14'd14839 : begin out <= 64'b0010010111000010101010001011001000101011000110101010000110001101; end
            14'd14840 : begin out <= 64'b1010101011101001001000110111110110101010011100010010101101010110; end
            14'd14841 : begin out <= 64'b0010101001010111000111011001100010011110010010001010011110111011; end
            14'd14842 : begin out <= 64'b0010100110000100100111111011100010101000100000101010101010011011; end
            14'd14843 : begin out <= 64'b1001100001101011101010101001111010101011101001001010010001111001; end
            14'd14844 : begin out <= 64'b1010100100101001101000011010111110100100101110001010011001010110; end
            14'd14845 : begin out <= 64'b1010101100010010100110001010111000100100100111100010101001001000; end
            14'd14846 : begin out <= 64'b1010010100111110001010101010100000011110001001001001110000110101; end
            14'd14847 : begin out <= 64'b1010100010001111001011000001000100101100001001100010101001001010; end
            14'd14848 : begin out <= 64'b1010100111110111001001101000111010101000111100110010100110101111; end
            14'd14849 : begin out <= 64'b0001010010100111001010001000101110101010000011111010100100111111; end
            14'd14850 : begin out <= 64'b0010000011010010101010110010111100101000101110000010100111000111; end
            14'd14851 : begin out <= 64'b0010101000001011101010100000010110101010000001010001111110111010; end
            14'd14852 : begin out <= 64'b0010011010110001101010100100110100100111111000001010101011011111; end
            14'd14853 : begin out <= 64'b0010011101110010101001101001001000101010101000000010010101010101; end
            14'd14854 : begin out <= 64'b1000100010100111001010100110111100100110000111010010010011001110; end
            14'd14855 : begin out <= 64'b1001011010011001001001100100101010101010000111000001100111111010; end
            14'd14856 : begin out <= 64'b1010011001000111101001101001101000100111101100011010100110111010; end
            14'd14857 : begin out <= 64'b0010001100101010101010011000000110101011011001010010100000011110; end
            14'd14858 : begin out <= 64'b1010000000101000101010101011110100011101001110110010101101111101; end
            14'd14859 : begin out <= 64'b1010101010001101101010111110110000101001100110000001111111001101; end
            14'd14860 : begin out <= 64'b1010010101100100001001001110110110101000111101111010100100110001; end
            14'd14861 : begin out <= 64'b1010101011111000101001001000001000101010010101111010100110010011; end
            14'd14862 : begin out <= 64'b0010010011010100101010010011010000101011001000101010010010101111; end
            14'd14863 : begin out <= 64'b0010100100100110101000010000100110100101111111001010101100001100; end
            14'd14864 : begin out <= 64'b1010010110111111101010111011100110011010111111010010101100100010; end
            14'd14865 : begin out <= 64'b0010101100101100001010111110010100011110111010100010011011011110; end
            14'd14866 : begin out <= 64'b1010010000100011001010101001010110101001011111101010101010000001; end
            14'd14867 : begin out <= 64'b0010101101100110101000110011111000011100010110100010010011001101; end
            14'd14868 : begin out <= 64'b1010100101010101101001101100011110100101000001011010011100100111; end
            14'd14869 : begin out <= 64'b0010010100000110001010100001010110101011010100100010100011000010; end
            14'd14870 : begin out <= 64'b0010101010101110001001100011000010101011011010010010000110101101; end
            14'd14871 : begin out <= 64'b0010000111100010101010111001110010011111111110111010010000010100; end
            14'd14872 : begin out <= 64'b1010001011100110101010101010010100101000010101000010011000001110; end
            14'd14873 : begin out <= 64'b1010010001100001001001100010111010101010101001101010101010010100; end
            14'd14874 : begin out <= 64'b1001111101001011001010001100110000100100101101111010001101111011; end
            14'd14875 : begin out <= 64'b1001100011101111101001010010101000101010010111010010101011000011; end
            14'd14876 : begin out <= 64'b0010011110010111001001000001010100011101011001100010011110101100; end
            14'd14877 : begin out <= 64'b0010001110010011000110111010001100101001011111011010011001001011; end
            14'd14878 : begin out <= 64'b0010101000001000000100010101100100011011100110011010001110000001; end
            14'd14879 : begin out <= 64'b0010100110001100001001001001101000100111110100001010011100010110; end
            14'd14880 : begin out <= 64'b0010010100000101001010100100000010101011011111010010101100110010; end
            14'd14881 : begin out <= 64'b1001101000101011100100111111000010101010011010101010101111111011; end
            14'd14882 : begin out <= 64'b0010001100110001101010100100101110101011011110011010101010001001; end
            14'd14883 : begin out <= 64'b1010100110110001100110100100011000011110110110111010101010101111; end
            14'd14884 : begin out <= 64'b1010010111000110001001100011010100100101011110011010101001011000; end
            14'd14885 : begin out <= 64'b1010101110110100101010000111010110011101101001010010100100011100; end
            14'd14886 : begin out <= 64'b1010101011101000000111010010110010101011000101111010001110100010; end
            14'd14887 : begin out <= 64'b0010000000100110000111111010101100100101001001111001110001111011; end
            14'd14888 : begin out <= 64'b1010100000000000001001110101001000100011000001001010100100001111; end
            14'd14889 : begin out <= 64'b1010101110100010001001111101110000011111111000101010000101101000; end
            14'd14890 : begin out <= 64'b1010101101101101101010111011001100010101011001011010100110000001; end
            14'd14891 : begin out <= 64'b0010011100001100001001110000010100100101100010011010100101011000; end
            14'd14892 : begin out <= 64'b0010010011001110101010010001101000101001100110100010100101000000; end
            14'd14893 : begin out <= 64'b1010101001010000001010011010010110100010001100101010011011000000; end
            14'd14894 : begin out <= 64'b0010101001110000101001100101010110100111001100110010100111100100; end
            14'd14895 : begin out <= 64'b1010101010110101101010010101110110100110001100101010011010011000; end
            14'd14896 : begin out <= 64'b1010001101011011100111110100010000101000110011000001000011111110; end
            14'd14897 : begin out <= 64'b1010000110111101101001110011110010100001000000100010000101001010; end
            14'd14898 : begin out <= 64'b0010011010111111101010000010110010100010011010010010010001110101; end
            14'd14899 : begin out <= 64'b1010010111100000101010011100111100101001101001011010001011111010; end
            14'd14900 : begin out <= 64'b0010000110100110101010011011111000100111110101000010000011100010; end
            14'd14901 : begin out <= 64'b0010100110110100101001101000000100100110110001111010100100101001; end
            14'd14902 : begin out <= 64'b0010001000010110101010110110110010101011100100111010000001011100; end
            14'd14903 : begin out <= 64'b1010100110101000101010001010101110100100000001010010000001100101; end
            14'd14904 : begin out <= 64'b0010100100111100001010111111000100101011000110101010101100101110; end
            14'd14905 : begin out <= 64'b0010100001011100000110001111010100100101100000100010100110000101; end
            14'd14906 : begin out <= 64'b1010100010111111101010110110110110101001100001001010101010110110; end
            14'd14907 : begin out <= 64'b1010101100010110001010001010100010011110010101110010011001110001; end
            14'd14908 : begin out <= 64'b1010011100001000001000100101011100011111001110110010101011001100; end
            14'd14909 : begin out <= 64'b1001111000100001101010010110101100101001110100001010010000000100; end
            14'd14910 : begin out <= 64'b1010100111000111001011000001011010101010010000010010011011010111; end
            14'd14911 : begin out <= 64'b0010100111100010001000101011011010100011010100010010001001000001; end
            14'd14912 : begin out <= 64'b1000010111101001101010001001110000101000111001111010101011101010; end
            14'd14913 : begin out <= 64'b0010010101010001101001010001111100101010001000010010100101101011; end
            14'd14914 : begin out <= 64'b0001100001001111101010011100111110101010100010011010011010101100; end
            14'd14915 : begin out <= 64'b0001111000111110100111111000010000100100001010010010011110111001; end
            14'd14916 : begin out <= 64'b1010011011101100001001010000101100100101100111001001111001100010; end
            14'd14917 : begin out <= 64'b0010000001000110001001011010101110101010011110001010010000010111; end
            14'd14918 : begin out <= 64'b0010000101010000101010101100010100101001111011011010011011011111; end
            14'd14919 : begin out <= 64'b1001100011110100101000001111011110101011110000101010011100000011; end
            14'd14920 : begin out <= 64'b1010100101111011101001000111011100100100110100000010011001011000; end
            14'd14921 : begin out <= 64'b0010101100001100101010101001100000101000000000001010100000100010; end
            14'd14922 : begin out <= 64'b0010011000111110001010001100011010100110001011101010101001101110; end
            14'd14923 : begin out <= 64'b1010000101000001001001010101001010101001000010110010100000011011; end
            14'd14924 : begin out <= 64'b1010010101100011000111000110111100100000100111000010011011101111; end
            14'd14925 : begin out <= 64'b0010000001010100001010001101101000100101010011001001110110101001; end
            14'd14926 : begin out <= 64'b1010010110111100101010011110110100100010011100111010100111111111; end
            14'd14927 : begin out <= 64'b1010101111110111101010000100001000100100111101001010101100111001; end
            14'd14928 : begin out <= 64'b0010101011001100001001010010101110100001101011011010100000000110; end
            14'd14929 : begin out <= 64'b0010100111110111101010010101001100011110010000011010101010100101; end
            14'd14930 : begin out <= 64'b0010010110000001001001100000100010101011010000011010001101101001; end
            14'd14931 : begin out <= 64'b1000110111010011001001010000110000101010000100110010000110111110; end
            14'd14932 : begin out <= 64'b0010010011100101101000010110111000011010001000110010100001001110; end
            14'd14933 : begin out <= 64'b0010010000101011100111010011110000100110010001000010100010101001; end
            14'd14934 : begin out <= 64'b0010101101100101101001111010100000101001100000010010101100101000; end
            14'd14935 : begin out <= 64'b1010010100011000001010001100111110101000111110001010101111000010; end
            14'd14936 : begin out <= 64'b1010101011011111000111101000101000100000000111010010100001110110; end
            14'd14937 : begin out <= 64'b1001110110100010101001101011001010100111110101110010101010110000; end
            14'd14938 : begin out <= 64'b1010000110101001101010010101101110101010011000100010101111010111; end
            14'd14939 : begin out <= 64'b1010101111101111101010001001000010100100110111001010100111101011; end
            14'd14940 : begin out <= 64'b0010110001011100101001111011110100100111101000111010100100011100; end
            14'd14941 : begin out <= 64'b1010101100111101100111110100101110101010011110001010101111111100; end
            14'd14942 : begin out <= 64'b1010101101110100101001100111000100100111101111100010001010110010; end
            14'd14943 : begin out <= 64'b0010011110000100001010100000110110101010000001010010101100011010; end
            14'd14944 : begin out <= 64'b1001100000001010001001011100111000101010110000001010011101010110; end
            14'd14945 : begin out <= 64'b1010101101011000101001110110101100101010011000000010100110100001; end
            14'd14946 : begin out <= 64'b1010000101100110101001001101001010100101000111100010100011111110; end
            14'd14947 : begin out <= 64'b1010101001110010001010010111100110101011011000100010010010101100; end
            14'd14948 : begin out <= 64'b1010100011011100001010110010100000101010000111110010010100111100; end
            14'd14949 : begin out <= 64'b1001111111010001001010111101010110100101010011111010000110111110; end
            14'd14950 : begin out <= 64'b1010100010001001001010010100110110101011011000101010100000010001; end
            14'd14951 : begin out <= 64'b0010100001011001001001110010000010101011101011001010101010010110; end
            14'd14952 : begin out <= 64'b0010011010010010101001000010000100011001100001101010100001101010; end
            14'd14953 : begin out <= 64'b0010101111011010101010010011100010100010011011100010101110100001; end
            14'd14954 : begin out <= 64'b1010101100100101101010010100010100100101010101011010011100111001; end
            14'd14955 : begin out <= 64'b1010011000001101101010100001000100100111100011010010001110100101; end
            14'd14956 : begin out <= 64'b1010100100010010101010000100101000100001101101011010010011010001; end
            14'd14957 : begin out <= 64'b1010101001100111001010100111011010100110100000000010011011101000; end
            14'd14958 : begin out <= 64'b0010100111100000001010010100010100100110010101110010010010000000; end
            14'd14959 : begin out <= 64'b1010010110000011101001110010000010100011111101100010101100111111; end
            14'd14960 : begin out <= 64'b0001101000101001101010000111111010101001001011010010010011000100; end
            14'd14961 : begin out <= 64'b1010010100111000001010101100111010101011001101111010100100110011; end
            14'd14962 : begin out <= 64'b0010100000100100001000011010101000100001000000000010011001111111; end
            14'd14963 : begin out <= 64'b1010100101011011101000010100111000101001110011111010011001101110; end
            14'd14964 : begin out <= 64'b0001100001000111001010110011110000101011000000111010100110000010; end
            14'd14965 : begin out <= 64'b0010100000101111101001110111001000101001011101111001110111010111; end
            14'd14966 : begin out <= 64'b1001011000010010001010011110000000101001110011111010100010110000; end
            14'd14967 : begin out <= 64'b0010100110101000001001100101000100101011011001000010101011111111; end
            14'd14968 : begin out <= 64'b0010001110010001101001011010010110101000001010110010100110100010; end
            14'd14969 : begin out <= 64'b0010101101111000001010101100101110101011100011011001111010100000; end
            14'd14970 : begin out <= 64'b1010010101011111000111010011110100101011110010000010101011111010; end
            14'd14971 : begin out <= 64'b1010010100101100101010011001011010101001110100011010101101010110; end
            14'd14972 : begin out <= 64'b1010011100101111101000011101011010101010001001001010100000111001; end
            14'd14973 : begin out <= 64'b1010100110000111101010111010100000101000000011010010100001010110; end
            14'd14974 : begin out <= 64'b0000111011110010001010011001110100101010010110001010001011100010; end
            14'd14975 : begin out <= 64'b0010011010000001001010101000110010101000110100000001111100010001; end
            14'd14976 : begin out <= 64'b0010011111001100100111110101000110100110011010100010001110011001; end
            14'd14977 : begin out <= 64'b0010100111110110001001011001111100011101000100001010100001101000; end
            14'd14978 : begin out <= 64'b1010010011101000001000100110010010100111101111010010010010110010; end
            14'd14979 : begin out <= 64'b0010000100010011101001000101111110101011001000001010101001001001; end
            14'd14980 : begin out <= 64'b1010010011111011101010110110100100100101101101011010101111001011; end
            14'd14981 : begin out <= 64'b0010101001001010000110101001000010100010001001100010110000010111; end
            14'd14982 : begin out <= 64'b0010011100101100000110111110010110100100000001001010011110100001; end
            14'd14983 : begin out <= 64'b0010011000100001001010010001111100100111010110101000110111011001; end
            14'd14984 : begin out <= 64'b1001100100001010001010100110001000011111010110011010101010111011; end
            14'd14985 : begin out <= 64'b0010010011100011101010101001000110100000101100011010100011000011; end
            14'd14986 : begin out <= 64'b0010010010111010101001010110111100010010001010001010101100111011; end
            14'd14987 : begin out <= 64'b0010001000010110001010011110110100100111001010000010011110100111; end
            14'd14988 : begin out <= 64'b0010101101000101101010011010000110101000010111010010101010010101; end
            14'd14989 : begin out <= 64'b1010011110000011001010110001100110101001110001111010101000100001; end
            14'd14990 : begin out <= 64'b0010010011000011101010101100001000011111111010000010001101100011; end
            14'd14991 : begin out <= 64'b1001110110110100101001010100110010101001111110100001111111111100; end
            14'd14992 : begin out <= 64'b0010010011001001101010010010011010011101100110010010100101011101; end
            14'd14993 : begin out <= 64'b0001011100110000001010111100100100101001100111110010101000010000; end
            14'd14994 : begin out <= 64'b0010101001010010001010100111001010001101110011110010101110110101; end
            14'd14995 : begin out <= 64'b0010101011100001101001000011110010100111100010110010101100111011; end
            14'd14996 : begin out <= 64'b0010100010000010101001111100111100101001101011101010100100101010; end
            14'd14997 : begin out <= 64'b0010000101110101100101101011010110101001000000101010001001011010; end
            14'd14998 : begin out <= 64'b0010100001110110001010100100000010101011011000110010010001001000; end
            14'd14999 : begin out <= 64'b1001100101001000101010011001100000011011010111010010101011001000; end
            14'd15000 : begin out <= 64'b1010010011101100001010101000111100101001000011011000001100111001; end
            14'd15001 : begin out <= 64'b1010000011010010001001100011010110100100011100011010101100110011; end
            14'd15002 : begin out <= 64'b1010100100011100001001011111010110101011101101110010101100011111; end
            14'd15003 : begin out <= 64'b0010101001000011001001011000011100101001101110101010101001111101; end
            14'd15004 : begin out <= 64'b0010100101101000101010100100010110100011000101011010000100011110; end
            14'd15005 : begin out <= 64'b0010000010000001001000010110011010101011100100011010101110010010; end
            14'd15006 : begin out <= 64'b0010100001000000101010100100101100100011100100010010100000110010; end
            14'd15007 : begin out <= 64'b1010100111011001101010100001100000100111111101111010011110101001; end
            14'd15008 : begin out <= 64'b1001010101011010001001100011011100101011101111100010101010011101; end
            14'd15009 : begin out <= 64'b1010011000110000101010101111100110101010101011100010101101111000; end
            14'd15010 : begin out <= 64'b1010101001001111101010011100111100100000000101011010000110110001; end
            14'd15011 : begin out <= 64'b0010001101101010001010111010100010100110110001000001100010111101; end
            14'd15012 : begin out <= 64'b0010101010011001001010110111001000100001000011000010100001000001; end
            14'd15013 : begin out <= 64'b1010101001101011101000010100101110101001001101001010101010110001; end
            14'd15014 : begin out <= 64'b0010010010001011001000101011111000011101001110101010011000110110; end
            14'd15015 : begin out <= 64'b1010100001011001001010000001101000101001010000011010011110001110; end
            14'd15016 : begin out <= 64'b1010000011000001100111000100010010010001111101110010011010001110; end
            14'd15017 : begin out <= 64'b1010100100001010101010110111111100100000011011001010100110000011; end
            14'd15018 : begin out <= 64'b0010101111010011001000101010101100101000011100110010011110010011; end
            14'd15019 : begin out <= 64'b0010000000100101101010011010001100011101110010001010000011101101; end
            14'd15020 : begin out <= 64'b0010101111110000001001001011001110011001110000111010100100011101; end
            14'd15021 : begin out <= 64'b1010010001100000101001101110011110100101001000111010101010010111; end
            14'd15022 : begin out <= 64'b1010101001101000101000101110011000101001001100111010001101110010; end
            14'd15023 : begin out <= 64'b1010100001010111001010100111001100101001011101001001111110000110; end
            14'd15024 : begin out <= 64'b1010010010101011101010011110010010100110110011110010100011110100; end
            14'd15025 : begin out <= 64'b0010101100010111001010000001010100100101010010011001110010000111; end
            14'd15026 : begin out <= 64'b0010100101001010101010110101111010001001001011000010011100101100; end
            14'd15027 : begin out <= 64'b1010011101111000001010011110010110101000000100111010011011100110; end
            14'd15028 : begin out <= 64'b0000111011100001101001111000100100101011001010010010100011111100; end
            14'd15029 : begin out <= 64'b0010101110000100001010000000101010101010000001101010100011000101; end
            14'd15030 : begin out <= 64'b0010101001110000101010000000011110011110101011001010101101111111; end
            14'd15031 : begin out <= 64'b1010101010111000000111110111001000011011100000110010101110110000; end
            14'd15032 : begin out <= 64'b1010010000110000100111110000100110101000010111001010000001101100; end
            14'd15033 : begin out <= 64'b0010101000110101001001101010011010101010000011010010100010100010; end
            14'd15034 : begin out <= 64'b0010010111000011101001000100100100101011000100101010100101011101; end
            14'd15035 : begin out <= 64'b0001001111010010101010101001111100101001100101111010011011010011; end
            14'd15036 : begin out <= 64'b1010010000111110101010001001110110000011000011100010100100100000; end
            14'd15037 : begin out <= 64'b1010100110000000101001011011001000100011010101011010000110100101; end
            14'd15038 : begin out <= 64'b1010101001010100101010000010000010011010101110001001110011111110; end
            14'd15039 : begin out <= 64'b0010101111001010101010101000111000101010100011010010011000001101; end
            14'd15040 : begin out <= 64'b1010010000000100001010100001110100010111000100000010100111000001; end
            14'd15041 : begin out <= 64'b0010000001110010001001110101100010101000101000000010101000010001; end
            14'd15042 : begin out <= 64'b1010010101000010101010001100110010100010101110110010101111111110; end
            14'd15043 : begin out <= 64'b1010010010010010001001001110111110100100100100111010011100010010; end
            14'd15044 : begin out <= 64'b1010100010111110001000000000110000101010001010110010101010101101; end
            14'd15045 : begin out <= 64'b1010000111100000101010000000110000100010100111101010101000111110; end
            14'd15046 : begin out <= 64'b1010000110010100001010101001111010100101011100100010011011010100; end
            14'd15047 : begin out <= 64'b0001110000110011101010010010110000100111000011110010100110100011; end
            14'd15048 : begin out <= 64'b1010101110111110101010000111001000101000100101101010101010010100; end
            14'd15049 : begin out <= 64'b1001111111001100001000000100101010101001011010000001111111110100; end
            14'd15050 : begin out <= 64'b1010101110111101001010110001011010100001101111001010100000111001; end
            14'd15051 : begin out <= 64'b0010101010000101101010000011011100101011110000010010101111110011; end
            14'd15052 : begin out <= 64'b1010110000011110001010110011101010101010000101110010010110110010; end
            14'd15053 : begin out <= 64'b0010101110101100101010010010001110100110111101001010010111111011; end
            14'd15054 : begin out <= 64'b1010100010010100101010111111000000010100000101110010100101111110; end
            14'd15055 : begin out <= 64'b0010101000011110101010011110100100100110110001000010011010001000; end
            14'd15056 : begin out <= 64'b0010101111100011001001011000101110100101101001110010100111101110; end
            14'd15057 : begin out <= 64'b1001110110101110100100010010010000100010010101000010100100010010; end
            14'd15058 : begin out <= 64'b0010001101010001001001001000110010101001001101010010100111100111; end
            14'd15059 : begin out <= 64'b1010101100011010001001001010011000101001110111100010100011101111; end
            14'd15060 : begin out <= 64'b0010101001110101001010110110001000101000101110001010100111001011; end
            14'd15061 : begin out <= 64'b1010100110011110101010110011110110101010000010100010010111101110; end
            14'd15062 : begin out <= 64'b1010101011100001001010010100110110100000000100100010100000101111; end
            14'd15063 : begin out <= 64'b0010101101000111001010010001100100101011001011101010100111110000; end
            14'd15064 : begin out <= 64'b0010100000000110100111111100001000101010100110111010011011100100; end
            14'd15065 : begin out <= 64'b0010101111101000000011100010001100101011000000001010101011110111; end
            14'd15066 : begin out <= 64'b1001100101100111001001100111101100100001111001101010100101110101; end
            14'd15067 : begin out <= 64'b1010100011000111100111011110100110100111010011011010101110110011; end
            14'd15068 : begin out <= 64'b0010101111100011001010011010001010100110000010101001111100010100; end
            14'd15069 : begin out <= 64'b1010011000110000001001110010010110101001100111011010100100001000; end
            14'd15070 : begin out <= 64'b1001111000011010000111000010000100101011101110101010100011011111; end
            14'd15071 : begin out <= 64'b1010010010110010001010011111001100101011100011010010100100001010; end
            14'd15072 : begin out <= 64'b0010001100010001001010100101101000100000100010100010100010101010; end
            14'd15073 : begin out <= 64'b0010100111000000000110011000101110101000000011110010010111101100; end
            14'd15074 : begin out <= 64'b1010011111111111100111110101000100001011111010100010101111011001; end
            14'd15075 : begin out <= 64'b1010101010001000001010111010000110101000001011011010000100011101; end
            14'd15076 : begin out <= 64'b0001000010010101101001110110110000101001111001001010000110100000; end
            14'd15077 : begin out <= 64'b0001110001101101001010101100010110100011010111000010011101000011; end
            14'd15078 : begin out <= 64'b1010101001101000101001010110010110100110111110100010000110100111; end
            14'd15079 : begin out <= 64'b0010110000111100001010011000001010101000110000110010011111110110; end
            14'd15080 : begin out <= 64'b1010000111111101001001100010000000100011110001110010010110101101; end
            14'd15081 : begin out <= 64'b0010011100001001101010101001001000101000011000100010100000100111; end
            14'd15082 : begin out <= 64'b1010100101110100101010011011011110100010101011101010110000000100; end
            14'd15083 : begin out <= 64'b0010010110001011001010010010110110101010011110001010101001001111; end
            14'd15084 : begin out <= 64'b1010010001001001101001111000110010101001100011101010011001011111; end
            14'd15085 : begin out <= 64'b0010011101110101001010001000100100100000100001000010101010110101; end
            14'd15086 : begin out <= 64'b1010001111001110001001110010100110100111110111001010100000001001; end
            14'd15087 : begin out <= 64'b0010000110110100101000011001100010101011000001001010100110111001; end
            14'd15088 : begin out <= 64'b0010100010110111001010011101101000100111101010010010001111010000; end
            14'd15089 : begin out <= 64'b0010001011000000101000101011111010100000100110100010100100001100; end
            14'd15090 : begin out <= 64'b1010011011000001000110111010100100101011100001100010010111000001; end
            14'd15091 : begin out <= 64'b1010101001110010100101101110100010101011001011001010100011010101; end
            14'd15092 : begin out <= 64'b1010000000110101001010100111010010101010011111101010100010110101; end
            14'd15093 : begin out <= 64'b0010000001100101100110110101101100101000001111110010101001001110; end
            14'd15094 : begin out <= 64'b0010100000011001001010010111111010101000111001110010011111110010; end
            14'd15095 : begin out <= 64'b1010101100101000101000110011111110011101011101011010101011010111; end
            14'd15096 : begin out <= 64'b1010011000011101101000101001110100101001110101001001111110100111; end
            14'd15097 : begin out <= 64'b0010101000101001101010100111101100101010010111000010010001000101; end
            14'd15098 : begin out <= 64'b0001100100110000101001101110001010101001000011000010100000011010; end
            14'd15099 : begin out <= 64'b0010101100011110101010110111001100100110001000011001110100100000; end
            14'd15100 : begin out <= 64'b0001111110100110001010100111111010100101111110100010010101110110; end
            14'd15101 : begin out <= 64'b1010101101110010101001111101100010100101010111100010010001011011; end
            14'd15102 : begin out <= 64'b1010010011010000001010011010001010100000011100001010010110010101; end
            14'd15103 : begin out <= 64'b1010100001010010101010011000101010100110101011111010101010001000; end
            14'd15104 : begin out <= 64'b1010100011011110001010001100010000100000010110010010101001111101; end
            14'd15105 : begin out <= 64'b1010100100000010101001111101000000100111000110100010010100101110; end
            14'd15106 : begin out <= 64'b0001110111110011100100000111111000101001001011001010001111000010; end
            14'd15107 : begin out <= 64'b1010100100100110101010010110110010100100101000101001110101001111; end
            14'd15108 : begin out <= 64'b1010100110100101001001101010100000101000001011000010101011000011; end
            14'd15109 : begin out <= 64'b0010100101111011101001110111011110101000000111111010000111101111; end
            14'd15110 : begin out <= 64'b0010011011101000001010111001111110101000001110111010001000000010; end
            14'd15111 : begin out <= 64'b0010100010110100101010111100100010100011010100010010011101011000; end
            14'd15112 : begin out <= 64'b1010010100101011101010010010000100100100010101101010011000111000; end
            14'd15113 : begin out <= 64'b1010010100011000001010110000011110100110101111111010101110010101; end
            14'd15114 : begin out <= 64'b0010010110111011001010001010010010100111111010001010010101111100; end
            14'd15115 : begin out <= 64'b1010100101000110101001010111110110101000011101101010101010000110; end
            14'd15116 : begin out <= 64'b0010001111001111001010111010001100100101110111100010100111111101; end
            14'd15117 : begin out <= 64'b1010010010111101001001000110110000101001010011101010100101000100; end
            14'd15118 : begin out <= 64'b0010101010100000101001000110000000011111011000001010011100100000; end
            14'd15119 : begin out <= 64'b1010100100010001001010011001010100101011010010101010011011110010; end
            14'd15120 : begin out <= 64'b0010100000010001001001100110111100100011101000011010101101111010; end
            14'd15121 : begin out <= 64'b0001111001111110001001101011101000101001011110001010011101010101; end
            14'd15122 : begin out <= 64'b0010101011111100101001011111011100101010011101001010000111100111; end
            14'd15123 : begin out <= 64'b1010101000000111001010101101100110101000011000001010001101101110; end
            14'd15124 : begin out <= 64'b1001111011001001001001101100011000101011000010100010011111100001; end
            14'd15125 : begin out <= 64'b0010100100001111001010100010101010011101001100101010101110000010; end
            14'd15126 : begin out <= 64'b0001111010111111001010101010001100100110111000111010101001000001; end
            14'd15127 : begin out <= 64'b0010110000000101001001000101000100101010000001011010101101111101; end
            14'd15128 : begin out <= 64'b1001110001010001001001111011001100101011101101111010100110100101; end
            14'd15129 : begin out <= 64'b0001001011101001001001001100010000100011010001011010100011111011; end
            14'd15130 : begin out <= 64'b1010001110011110001010000111011100100001111101100010010101100110; end
            14'd15131 : begin out <= 64'b0010000000001011000111001111101110100110011110011010101101010010; end
            14'd15132 : begin out <= 64'b0010101100011101001010110001001110101011001111110010011010010101; end
            14'd15133 : begin out <= 64'b1010001011111110000110100100101100101000101011111010010110000111; end
            14'd15134 : begin out <= 64'b0010100011110011101010101101001110101010000101111010101111011111; end
            14'd15135 : begin out <= 64'b0001010111110010101010011010010110100110011010101010100111111001; end
            14'd15136 : begin out <= 64'b0010001110101011101001010110111010100111101111001010000100001010; end
            14'd15137 : begin out <= 64'b1010100010111111101010100110000010101000010001101010100001100011; end
            14'd15138 : begin out <= 64'b0010001010010111001010010101111000011011110100000010001000001000; end
            14'd15139 : begin out <= 64'b1010001001100100101010110101010100100111101001001010011100100110; end
            14'd15140 : begin out <= 64'b0010100011111001001010010011100110101010110110000010101000011001; end
            14'd15141 : begin out <= 64'b1010000110010100001010100101110010100001001111100010100111101101; end
            14'd15142 : begin out <= 64'b1010001000110011001001001111011010101000011001001010001010011111; end
            14'd15143 : begin out <= 64'b1001110001011111001010111100000010011101101010100010100010000010; end
            14'd15144 : begin out <= 64'b0010010001100001101010001010111100100101111010111010001000101100; end
            14'd15145 : begin out <= 64'b1010101110101100101010101000110100101001011001101010010100010101; end
            14'd15146 : begin out <= 64'b1010101100000001101010011001101100101001010011101001110000000101; end
            14'd15147 : begin out <= 64'b1010100000101110001010010101011000100111001010001010100101010000; end
            14'd15148 : begin out <= 64'b1010101001000001100111000101001110101011011110001010011101011000; end
            14'd15149 : begin out <= 64'b0010101000100111001010001111101110101010000111111001010001110111; end
            14'd15150 : begin out <= 64'b1001011101100010001010000111100100101000100011001010010000001010; end
            14'd15151 : begin out <= 64'b1010100000001000100110011111110000101010010010000010100101011111; end
            14'd15152 : begin out <= 64'b1010010011000101001001101110111000100000111001010010010101000100; end
            14'd15153 : begin out <= 64'b1010100101111010101001100101001100011001000010110010010110000100; end
            14'd15154 : begin out <= 64'b1010100111101110001010110011000110101000010110100010100011101101; end
            14'd15155 : begin out <= 64'b1010101000011111101010010111100110101011110011110010001111001100; end
            14'd15156 : begin out <= 64'b0010010110111000101010000110101100011100011101001010000010111000; end
            14'd15157 : begin out <= 64'b0010001110111110100110101100101000101011001111111010100110000110; end
            14'd15158 : begin out <= 64'b0010011010100100001010110101011000101001111111001010010110101111; end
            14'd15159 : begin out <= 64'b0010101101011010101001111101101000101010100010010001100011000000; end
            14'd15160 : begin out <= 64'b0010101111001001101010011110111010101011001001010010101111110101; end
            14'd15161 : begin out <= 64'b0010000000001001101000011010100000011101000110011010101000101110; end
            14'd15162 : begin out <= 64'b0010101101011101101010101010101110100111101101110010000110001100; end
            14'd15163 : begin out <= 64'b0010100111000000101001001011001100101001100101111010001011101101; end
            14'd15164 : begin out <= 64'b0010100111011001001010000110101100101000010011110010101011101000; end
            14'd15165 : begin out <= 64'b1010011101101011101010011000101000101011011110100010000100010110; end
            14'd15166 : begin out <= 64'b0001110110101110001010000110011010101010101100010010010001100010; end
            14'd15167 : begin out <= 64'b0000110100110011001001000000011100100011110101111010100110101110; end
            14'd15168 : begin out <= 64'b0010001000101010000110101011010010101001101000010010101111010000; end
            14'd15169 : begin out <= 64'b0010001111001011001011000011011010100100101110000010100101000001; end
            14'd15170 : begin out <= 64'b1010011001100001101010111101011110100110011101100010100010101001; end
            14'd15171 : begin out <= 64'b0000010100001110001001000010010110100110101101100010101111000101; end
            14'd15172 : begin out <= 64'b1010011100101000101001011100010010100010011010110001110001011111; end
            14'd15173 : begin out <= 64'b1010011100100001101010110010100110101000000111101010100011011010; end
            14'd15174 : begin out <= 64'b0010101000011001101001010110000010100000001100110010101001111110; end
            14'd15175 : begin out <= 64'b0001100110001101101010101101100000010100110010100010011000001111; end
            14'd15176 : begin out <= 64'b1010001001011101000111101110111010101000001001001001110110100001; end
            14'd15177 : begin out <= 64'b1010101100011011100111110110000100100101000010010010100001001010; end
            14'd15178 : begin out <= 64'b0010100011111000101001011000111000100110111111101001110011111101; end
            14'd15179 : begin out <= 64'b1010100110000011101010101011010010100000111011000010101010110001; end
            14'd15180 : begin out <= 64'b1010011000011010000111000100001110010101110100000010001100011110; end
            14'd15181 : begin out <= 64'b0010001100111111001001010110001000101010100110100010100000011011; end
            14'd15182 : begin out <= 64'b0010100000001111101010010001010010101000011000011010101001000011; end
            14'd15183 : begin out <= 64'b1010000001101101001001000100101100100001010010010010101111110001; end
            14'd15184 : begin out <= 64'b1010000111111011101010000001001000100111101100100010010100000101; end
            14'd15185 : begin out <= 64'b1010001011000111101000011011011110100110100000000010101001011111; end
            14'd15186 : begin out <= 64'b0010100010101100001010110010100000101011010101001010100010111101; end
            14'd15187 : begin out <= 64'b1010101100111100001001010001000100101010000010001010001011101100; end
            14'd15188 : begin out <= 64'b1010101101111001001010001011001010101010111101010010011111110100; end
            14'd15189 : begin out <= 64'b1010100110011001001010001111111010101011001100010010011011010010; end
            14'd15190 : begin out <= 64'b1010100100001011101000000101111010101000100111100010011001001100; end
            14'd15191 : begin out <= 64'b1001101110100010101010010101000010101001110101100010101111000010; end
            14'd15192 : begin out <= 64'b0001110010010110001001001111100110101010101111101010100000001000; end
            14'd15193 : begin out <= 64'b1010010010000100101000010010111110101000111100110010101110101010; end
            14'd15194 : begin out <= 64'b0010101000010000101000000110001000101010101110101010011011111000; end
            14'd15195 : begin out <= 64'b0001000100001101001010010101011100100101101110110010101111111111; end
            14'd15196 : begin out <= 64'b1010100010011010001010000110111010011000101100110010101101100001; end
            14'd15197 : begin out <= 64'b1010100000110011001000110000010110100101000011110010101111101000; end
            14'd15198 : begin out <= 64'b1001111111100101101010100101010110101010100011001010011101011100; end
            14'd15199 : begin out <= 64'b1010100001110110101001100000010000100010110010111010100010101101; end
            14'd15200 : begin out <= 64'b1010100001101000000111100101111010101011101011101010100010110111; end
            14'd15201 : begin out <= 64'b1001101001000100001010000101110110101001000101001010100100000111; end
            14'd15202 : begin out <= 64'b1010101100011111001010000010100110101011111001001001110001101111; end
            14'd15203 : begin out <= 64'b0010011001001101101000101101000110101011111101001010100110000101; end
            14'd15204 : begin out <= 64'b0001010101101001001010000100101010101001101100011010100111000000; end
            14'd15205 : begin out <= 64'b0010101001111110001010001010000010011110010000110010000101011100; end
            14'd15206 : begin out <= 64'b1010010101011000101001001001000010101011000011010010101110000101; end
            14'd15207 : begin out <= 64'b0010100100111101101001101111000100100111010000000010101100001000; end
            14'd15208 : begin out <= 64'b1010011011001110001001100110000000011001010100101010001011100001; end
            14'd15209 : begin out <= 64'b0010100011111000101000100100100010100010010101000010010000110111; end
            14'd15210 : begin out <= 64'b1010101100101000001001100100100100100001010001111001110111111110; end
            14'd15211 : begin out <= 64'b0010101001101110101000100111000000101001110100000010101011101001; end
            14'd15212 : begin out <= 64'b0010100101100011101010100011100110100111101000100010101101101101; end
            14'd15213 : begin out <= 64'b1010101001000001101010110000101010101010100100011010100000001001; end
            14'd15214 : begin out <= 64'b0010011111100110001001110010100110100100001010011010000100101010; end
            14'd15215 : begin out <= 64'b1010101001010011000111110101000100100101000010111010010000111101; end
            14'd15216 : begin out <= 64'b1010101001110010101010010011110000101010101000011010101111111110; end
            14'd15217 : begin out <= 64'b1001111100111000101010111011000000101011011000000010101010111100; end
            14'd15218 : begin out <= 64'b0010101111100011101001110010001100101011100001011010000111001101; end
            14'd15219 : begin out <= 64'b0010101100101101101010110110010010101010111100010010001100001000; end
            14'd15220 : begin out <= 64'b1010010000101010101001001110100000100100010010101010000111001100; end
            14'd15221 : begin out <= 64'b1010100011000100001001100100100100100110100100011010100111111010; end
            14'd15222 : begin out <= 64'b1010101111110011101010011100111110100111101010101010011001011101; end
            14'd15223 : begin out <= 64'b0010110001100110001001010001111100011111111001000001110001110001; end
            14'd15224 : begin out <= 64'b0010101010100100100110111001010110101010001001001010010011100011; end
            14'd15225 : begin out <= 64'b0010011010101100101001010000110010101000001010010001100000101101; end
            14'd15226 : begin out <= 64'b1010011110010101000110110100110010101001101001101010100000110101; end
            14'd15227 : begin out <= 64'b0010000010100100001010000111010000101001011000000010100010000000; end
            14'd15228 : begin out <= 64'b0001100110111101001010011101010000100011000001111010010101111000; end
            14'd15229 : begin out <= 64'b1001111000010100100110001001001000100100011000100010011000111111; end
            14'd15230 : begin out <= 64'b0001100110111110001001011100011000101000000101101010011100001000; end
            14'd15231 : begin out <= 64'b1010011111001110101010011011000010011000111001001010100100011101; end
            14'd15232 : begin out <= 64'b0010100101010101101010110011100100101000111110100010100101000011; end
            14'd15233 : begin out <= 64'b0010110000000001101000000011001000100010010111111000001000000010; end
            14'd15234 : begin out <= 64'b0010000011100111001010001101000100100001000101110010101111100010; end
            14'd15235 : begin out <= 64'b0010011101101000001001011110111010100111000111100010100100001001; end
            14'd15236 : begin out <= 64'b0010000100010000101000110111100010100010100100110010101000000001; end
            14'd15237 : begin out <= 64'b1001110000110010101010010010101100101010001110110010100000100100; end
            14'd15238 : begin out <= 64'b1001010100000100001010011100001000100000101010001001110010011001; end
            14'd15239 : begin out <= 64'b1010101110011111101010111110110000101000111011111010001001000110; end
            14'd15240 : begin out <= 64'b0010010001000100001010101010100100101001110011100010101000001011; end
            14'd15241 : begin out <= 64'b0010101100101010001000011001011000011001001111110010100101010111; end
            14'd15242 : begin out <= 64'b0001111110100001001010111111011100101011111100010010100100001111; end
            14'd15243 : begin out <= 64'b0010011111101101001001011001010000100010111101011010100110010110; end
            14'd15244 : begin out <= 64'b0010000010000010001001111001101110100010110011000010101111001001; end
            14'd15245 : begin out <= 64'b0010100110111110101010111000000110011000101000001010101101111101; end
            14'd15246 : begin out <= 64'b1001101111110100001001000111100010101011100101010010010000100100; end
            14'd15247 : begin out <= 64'b1010010001111011101010100011010000101010010011101010100111110011; end
            14'd15248 : begin out <= 64'b1010101001101010101010111111010000101010111000101010011011111010; end
            14'd15249 : begin out <= 64'b0010000010011110001010010011010010101010011001101010101001011011; end
            14'd15250 : begin out <= 64'b0010001010101011001010001001100110101000010001111010010000101000; end
            14'd15251 : begin out <= 64'b0010100110111001000111010010111100011010010110110010100110010110; end
            14'd15252 : begin out <= 64'b1010110000001110001010110001000010101000010011101010101011001100; end
            14'd15253 : begin out <= 64'b0000001101010011101001110111111000101011011010101010010010001011; end
            14'd15254 : begin out <= 64'b0010011100010111101010110100001000100110000100110010101101110000; end
            14'd15255 : begin out <= 64'b0010000010011100001010001010100110100100101001011010100001001110; end
            14'd15256 : begin out <= 64'b0010011010011100101010110011010100101000001110010001110010010101; end
            14'd15257 : begin out <= 64'b0010100110001010101001001101000100100111100110000001011100011100; end
            14'd15258 : begin out <= 64'b1010100101100000101001100011100010101001011000000010010010000001; end
            14'd15259 : begin out <= 64'b0010010000110101101010111111000010101011101001100010100000111101; end
            14'd15260 : begin out <= 64'b1010101110101011101010110001111010100011111101101010101001110011; end
            14'd15261 : begin out <= 64'b0010010110100110000111001011000000100111100101100001010111001110; end
            14'd15262 : begin out <= 64'b0010110000010001000101101110101010100001110100101010001100111111; end
            14'd15263 : begin out <= 64'b0010010101110101001010001001000010100110001011000010101011110101; end
            14'd15264 : begin out <= 64'b1010101011000001100111100111011000101000001001001010100000000100; end
            14'd15265 : begin out <= 64'b1010001101110011001001011100000110100010101010101010000100000010; end
            14'd15266 : begin out <= 64'b1010010000100101101010000100101010100011101001010001110010100101; end
            14'd15267 : begin out <= 64'b1010001110101110101011000100000100101000101011001010010100101101; end
            14'd15268 : begin out <= 64'b0010100011000000001001100010011010101011101110001001110100110001; end
            14'd15269 : begin out <= 64'b1010100101000101001000011001000010101000100000100010100010010101; end
            14'd15270 : begin out <= 64'b1010101110111111101001110101001100100100011010111010100100001101; end
            14'd15271 : begin out <= 64'b0001100110001011001001011011100010101001010110101010010101101101; end
            14'd15272 : begin out <= 64'b1010000111000010001000101110100100100010111001000001111100111111; end
            14'd15273 : begin out <= 64'b0010010011110110101010100010010100101000001000000010101011011100; end
            14'd15274 : begin out <= 64'b1010100101110110101000101111110010101011100000101010101111110000; end
            14'd15275 : begin out <= 64'b1010010100000001101010010001011010011101110101110010101011001110; end
            14'd15276 : begin out <= 64'b0010100100100000001010011000001110101001011001101001111100110111; end
            14'd15277 : begin out <= 64'b0010101101011011001010100110100100101011110101000010100110100001; end
            14'd15278 : begin out <= 64'b1010100001001111001001100101111010101011101010111010011000011011; end
            14'd15279 : begin out <= 64'b1010010010001111001000000111100100100101101111111010001001101001; end
            14'd15280 : begin out <= 64'b1010010010101100000111000101110010101000001111101010100001011000; end
            14'd15281 : begin out <= 64'b1010100011111100101010111001100110101010100000010010100101001100; end
            14'd15282 : begin out <= 64'b0010001100110010100111100111000110100011011111000010100101101101; end
            14'd15283 : begin out <= 64'b1010101101011011100011111000111100100010111100001010011100000101; end
            14'd15284 : begin out <= 64'b1010101011010111001010000010110100101000111011000000110110001111; end
            14'd15285 : begin out <= 64'b1010001001010100001010101000101100011101111111010010001000010010; end
            14'd15286 : begin out <= 64'b1010100111101111001010101101001110010010010011010010101010001011; end
            14'd15287 : begin out <= 64'b0010100000101001001001010111000010100000010110110001001000101000; end
            14'd15288 : begin out <= 64'b1001110111010011001000010110101100101000011101000010010010111001; end
            14'd15289 : begin out <= 64'b0010010010010101000111010111100000100110011000001010010001011100; end
            14'd15290 : begin out <= 64'b1010011101111111001001101010011100100111100101101010010110011110; end
            14'd15291 : begin out <= 64'b0010100011001111101010000000101010100111110111110010000110010000; end
            14'd15292 : begin out <= 64'b1010100000100111101010011110011110101011111110111001110010001000; end
            14'd15293 : begin out <= 64'b1010000000110110100110100101001010101000111010101010101001011100; end
            14'd15294 : begin out <= 64'b1010101001110101101010010000010010101001001000111010101111000110; end
            14'd15295 : begin out <= 64'b0001101110110010001000000111000100101011110010101010011110101101; end
            14'd15296 : begin out <= 64'b0010101011001010001011000000100000101010110011011001100011111001; end
            14'd15297 : begin out <= 64'b0010100100000010001010111010000100100100110111001010101010011101; end
            14'd15298 : begin out <= 64'b0001011000101110101001111110010110100001011111100010100110000111; end
            14'd15299 : begin out <= 64'b0010011100011101101001011110011000101010001011001010100000001011; end
            14'd15300 : begin out <= 64'b0000101101011100101000100001111110100111011011001010010111010010; end
            14'd15301 : begin out <= 64'b0010101110000101101010011110101010100110111000101010011001111101; end
            14'd15302 : begin out <= 64'b1010101111111010001010100010100110100101000100100010000010101111; end
            14'd15303 : begin out <= 64'b1010010101100110101010011101111100100111111110111010011000101110; end
            14'd15304 : begin out <= 64'b1010010110011111001010111111010010101000111101011010101111000101; end
            14'd15305 : begin out <= 64'b1010000010000001001010110101010010100111100101000001011110100101; end
            14'd15306 : begin out <= 64'b0010010000001010100111110110001010101001101010010001001000111001; end
            14'd15307 : begin out <= 64'b1001100100000010001000111011000000101000000111111010000100000111; end
            14'd15308 : begin out <= 64'b0001011100010101000111000011111010010011000100100010100110010011; end
            14'd15309 : begin out <= 64'b0010011101111010101010111000101000100100100100101010000011101111; end
            14'd15310 : begin out <= 64'b0010101110010000001001010100101000010100101110100010001110011100; end
            14'd15311 : begin out <= 64'b0010101000100010101000101100101110010101111010010010010010111010; end
            14'd15312 : begin out <= 64'b0010100001000000101000001000000010100010100010001010001010110100; end
            14'd15313 : begin out <= 64'b1010100111100001001010100100011000100011100110010010100010010010; end
            14'd15314 : begin out <= 64'b1001110011001001001000111101110010100101101101001010100011000011; end
            14'd15315 : begin out <= 64'b0001111011000110101010011000110110100001010111010010011001111010; end
            14'd15316 : begin out <= 64'b0010100000000111001000100001001100100101010000100010011110000111; end
            14'd15317 : begin out <= 64'b0010101101000111101010000100011010101000001100110010100011101001; end
            14'd15318 : begin out <= 64'b0001111000011000101001110101011000100101011101100010100110001100; end
            14'd15319 : begin out <= 64'b0010100000010111001010001000101110011101111100101010011000011100; end
            14'd15320 : begin out <= 64'b0010100010011111101001001011001110100111101001001010101101111000; end
            14'd15321 : begin out <= 64'b0010110001110000001010001010100010101010100000100001111100110111; end
            14'd15322 : begin out <= 64'b0010101000011010101010101000101100101010010010110010101000111010; end
            14'd15323 : begin out <= 64'b0010100110000101101010100011001010100101101011001001111001001000; end
            14'd15324 : begin out <= 64'b0010001110010111101010110010100110100110000111100010101111110110; end
            14'd15325 : begin out <= 64'b0001100110100111001010101100010110011101110100010010001010110101; end
            14'd15326 : begin out <= 64'b1010101101110111001010011010001010101011011101001010010111010100; end
            14'd15327 : begin out <= 64'b0010100010100010001001001101110110100100101000110001111001100111; end
            14'd15328 : begin out <= 64'b0010000001111010101010010011011110101011101010101001100101001011; end
            14'd15329 : begin out <= 64'b0010100011100011101000010111111010101000100011101010101011011101; end
            14'd15330 : begin out <= 64'b0010011100110101001010001000101010101001011010010010100011001011; end
            14'd15331 : begin out <= 64'b0010000010001100001001100000000110011100001001010010100011110100; end
            14'd15332 : begin out <= 64'b0010011101010010001001011010000000101010111100101001110100011111; end
            14'd15333 : begin out <= 64'b0010100001110010001010011010011010100100100011011010100110101010; end
            14'd15334 : begin out <= 64'b0010100111000111001010101101010010101010111010100010010111000011; end
            14'd15335 : begin out <= 64'b0001101100001011101010100011100000101010110110111010001111011111; end
            14'd15336 : begin out <= 64'b0010101100011111101010001011010000101001001001110010101111101000; end
            14'd15337 : begin out <= 64'b0010001101100101100111011100101000101001100111000010011100110000; end
            14'd15338 : begin out <= 64'b0000111100100000101010101110001110101011000100101010000100000010; end
            14'd15339 : begin out <= 64'b0001000000100100001000010110111110100001001101001010100110001101; end
            14'd15340 : begin out <= 64'b0010011000001111001010010101001110100010010100111010100011110101; end
            14'd15341 : begin out <= 64'b1010100111111000001000011001100100101011010111001010010101100000; end
            14'd15342 : begin out <= 64'b0010100100111000101010010000100110011110000100000010101101100111; end
            14'd15343 : begin out <= 64'b0001111011001010001001001101010100101011101111011010000000000001; end
            14'd15344 : begin out <= 64'b0010100100111010100111101010000110101010101011100001111111100100; end
            14'd15345 : begin out <= 64'b0001010111110100101001111001001010100111001001111010100011111001; end
            14'd15346 : begin out <= 64'b0010000001100010001010100010010110101010101010100010011100111011; end
            14'd15347 : begin out <= 64'b1010101011010000000100100011111100101011010110110010101010000011; end
            14'd15348 : begin out <= 64'b0010101101101101101010001100111010101001100000000010010111001011; end
            14'd15349 : begin out <= 64'b0001100100001101001010001110100110101011011110110010010010110011; end
            14'd15350 : begin out <= 64'b0010011011011001001010001011111110101001011111100010011011100011; end
            14'd15351 : begin out <= 64'b0010101110101000101001101001111010101001000001110010010011100010; end
            14'd15352 : begin out <= 64'b1010100100000111101010101111111010101010110010010010100100001100; end
            14'd15353 : begin out <= 64'b0010101100000011001001110110111000101000111001110010101000110001; end
            14'd15354 : begin out <= 64'b0010100010111000001010101010000100100010111110101001110111110001; end
            14'd15355 : begin out <= 64'b0010011000000001001001101010001010011111010010110001101111100011; end
            14'd15356 : begin out <= 64'b0010001100001100001000001101000100101011000010110010101100010110; end
            14'd15357 : begin out <= 64'b1010001001001101000111010001100100101011100001000010000001011111; end
            14'd15358 : begin out <= 64'b1010011011000011101000111011101000100111100111111001101000010010; end
            14'd15359 : begin out <= 64'b1010000100111010101000011101110110100110011100010010001010110001; end
            14'd15360 : begin out <= 64'b1010000000011011101001110001100110101001001001110010101000101110; end
            14'd15361 : begin out <= 64'b1010101100011100101000000110100000100111000110111010100000101101; end
            14'd15362 : begin out <= 64'b0010100100010101001010001010000100100101101111101010101001100100; end
            14'd15363 : begin out <= 64'b1010000010110110101010011100101010100101100110000010100011100010; end
            14'd15364 : begin out <= 64'b1010101100000101001010110110010010100111111011110001110000100011; end
            14'd15365 : begin out <= 64'b0010010011000111101010111010000000100001111010111010010110111011; end
            14'd15366 : begin out <= 64'b0010101111001010101010111011110010101010100100100010000010101001; end
            14'd15367 : begin out <= 64'b1010101000100101001010010101111000100000010010100010011100111110; end
            14'd15368 : begin out <= 64'b0001111011000001101010011001110010100100000000011001111101010101; end
            14'd15369 : begin out <= 64'b1010101110000101101010110000000110100101100010101010100001110010; end
            14'd15370 : begin out <= 64'b0010000101001111001001011110000010101000000000110010011001111001; end
            14'd15371 : begin out <= 64'b1010101010000010101010101011011110101000001100001010100001101010; end
            14'd15372 : begin out <= 64'b1010011001001111001000010100100000100111111111001001000110001001; end
            14'd15373 : begin out <= 64'b1010010011000011101001101101110000101010100011000010101101100110; end
            14'd15374 : begin out <= 64'b1010010111100000001010110100110000100100110110100010100010101010; end
            14'd15375 : begin out <= 64'b0010011110101100001010111001101100001010000010100010101001000010; end
            14'd15376 : begin out <= 64'b1010011000010101101010110100101000101001100001000010100011100001; end
            14'd15377 : begin out <= 64'b1010010000010000101010011100111000100011111011101010001110000001; end
            14'd15378 : begin out <= 64'b1010011011100101001010001110001110101001100110100010011010110101; end
            14'd15379 : begin out <= 64'b0010100011010000001010010000011110101000000001011010011111001001; end
            14'd15380 : begin out <= 64'b0010010010000010001001110001000100100011101010010010010101011100; end
            14'd15381 : begin out <= 64'b0010100011111010001010010010011000101010010011110001011001110000; end
            14'd15382 : begin out <= 64'b1010101000010101001010001110010010100111010000111010101111011001; end
            14'd15383 : begin out <= 64'b1010011010101001000111000110100110100100011111001010101000011111; end
            14'd15384 : begin out <= 64'b1010101001010110100110111011000010101011011010101010101010101011; end
            14'd15385 : begin out <= 64'b1010000110101010001001000100001010101001000000011010101101111100; end
            14'd15386 : begin out <= 64'b0010010011100001101010110110010010100110001000100010010110011010; end
            14'd15387 : begin out <= 64'b1010100110100111001010101100001010101000011011111010100000101000; end
            14'd15388 : begin out <= 64'b0010100110010010001010111101010100100101000101101010010001010110; end
            14'd15389 : begin out <= 64'b1010100100000001101010100010010000101001010101111010101000110011; end
            14'd15390 : begin out <= 64'b1010010100011110001011000110010100100101011110100010000101010110; end
            14'd15391 : begin out <= 64'b1010100000110100101010011111001100100101100101000010100111101111; end
            14'd15392 : begin out <= 64'b0010101001101110001001110011100100100111011000101010001101100101; end
            14'd15393 : begin out <= 64'b0010101000110010101010000001000000101011101010111010100101011111; end
            14'd15394 : begin out <= 64'b0010010101100111101001111010001110101001010000101010101001101001; end
            14'd15395 : begin out <= 64'b1010011110011000001001010111000010101010001111000010010001101010; end
            14'd15396 : begin out <= 64'b0010011111011100000110000001000010101000101100110010100100110110; end
            14'd15397 : begin out <= 64'b1010101100000011101000011100011100101000111001110001111010101011; end
            14'd15398 : begin out <= 64'b0010100010001100101010010001101000100001110101000010101110100000; end
            14'd15399 : begin out <= 64'b1010101111101010000011000000010100100100011111001010010010101010; end
            14'd15400 : begin out <= 64'b1010100001001100101001000011100010100011011101001010101001000001; end
            14'd15401 : begin out <= 64'b1010011010101111001001100110110000101000111101100010101010100111; end
            14'd15402 : begin out <= 64'b1010001110111010001000010101011110101001100110110010010101010010; end
            14'd15403 : begin out <= 64'b1010011001110000001010001100111110101010111000100010011101111000; end
            14'd15404 : begin out <= 64'b1010100110100111001010001001111000100100000101101010011001101010; end
            14'd15405 : begin out <= 64'b0001110100101011001001010011011110101011111110001001111111101010; end
            14'd15406 : begin out <= 64'b0010011110000110101001100010100110100110110011000001110011010111; end
            14'd15407 : begin out <= 64'b1010010111101111001001010111111010100110010000101010101100010010; end
            14'd15408 : begin out <= 64'b1010010101001111001010100111100000100110111011101010101111101111; end
            14'd15409 : begin out <= 64'b0010100011010111101001001010111110101000101001111010101101001111; end
            14'd15410 : begin out <= 64'b1001110111110111001010110011100010101011011110000010101011110000; end
            14'd15411 : begin out <= 64'b0010101100111010001010011010001000101010001010100010011010001101; end
            14'd15412 : begin out <= 64'b1010011101110001001000010011110010100111110011101010010001101101; end
            14'd15413 : begin out <= 64'b1010101101000111001010001110101110100111010011100010100001000110; end
            14'd15414 : begin out <= 64'b1010001111000100001010000001100110101000010000101010101011010111; end
            14'd15415 : begin out <= 64'b1010101110101110001001000111110010100000100010110010100110000001; end
            14'd15416 : begin out <= 64'b1010010100011111101010100111010100100101110111000001001100000101; end
            14'd15417 : begin out <= 64'b0010010010101111001010010010111100101001111010110010100011000000; end
            14'd15418 : begin out <= 64'b0010101100001110101010000011100010101000110101000010100100101100; end
            14'd15419 : begin out <= 64'b0010100111010000101001010110101010100100011000100010101010110111; end
            14'd15420 : begin out <= 64'b0010100010101010001010001011111010100001011000101010010010110111; end
            14'd15421 : begin out <= 64'b0010010000011110001000100110010000101011001101010010101010101000; end
            14'd15422 : begin out <= 64'b0010100011100011001001111101001000100110110111111010100101111010; end
            14'd15423 : begin out <= 64'b0001110100101100001001100101100110100100011101010010011110100010; end
            14'd15424 : begin out <= 64'b1001111100011100001001100100110010101000011010001010101111100001; end
            14'd15425 : begin out <= 64'b1010100001000000101001010010110010100110000110100010101010000100; end
            14'd15426 : begin out <= 64'b1010011011000110101010101011001010101001001111110010010001011000; end
            14'd15427 : begin out <= 64'b1010100001111000001010110110001100100000001000011010101100100000; end
            14'd15428 : begin out <= 64'b1010100010001010001010110011000010100100000010100010101111000111; end
            14'd15429 : begin out <= 64'b0010101000100101001010101000111100101001110010110010100001110101; end
            14'd15430 : begin out <= 64'b0010101111111101001010001101100000100110010101011010100100100100; end
            14'd15431 : begin out <= 64'b1010110000000000101010000011000100101001110010111010100011100000; end
            14'd15432 : begin out <= 64'b0010001011101110001010101000011000101000111000110010011010111101; end
            14'd15433 : begin out <= 64'b1010101100000001000111010100110000101001101001100001101001000100; end
            14'd15434 : begin out <= 64'b1010101100000100001000001100000110101001101000100010100001111000; end
            14'd15435 : begin out <= 64'b1010101010100011101010100111001100010101111011100010100000110011; end
            14'd15436 : begin out <= 64'b0010100000010000001010100011001110100101001001001010000011001011; end
            14'd15437 : begin out <= 64'b1010011001000011101000010010100000100100000110101010100011101101; end
            14'd15438 : begin out <= 64'b1010010101110011001010000110111100100111111100101010100111100110; end
            14'd15439 : begin out <= 64'b1010010010000111001000110101011100101001111111011010010001000110; end
            14'd15440 : begin out <= 64'b0010000000011000101010110100001100101001010001001010100101101100; end
            14'd15441 : begin out <= 64'b0010100011100001101011000001100000011000000111100010100000010001; end
            14'd15442 : begin out <= 64'b0010101001000011101010001101111110101011100111001010100011110000; end
            14'd15443 : begin out <= 64'b0010011010111010100111010011001000100010110000010010100110010000; end
            14'd15444 : begin out <= 64'b0010101001110100101010000111001100101010101001000010100001111010; end
            14'd15445 : begin out <= 64'b0010101100011001001001111010010100101000010011011010001111110001; end
            14'd15446 : begin out <= 64'b0000110101100011101001011100000000101100000101110010001110100011; end
            14'd15447 : begin out <= 64'b0010001100011011001010000011111000101001111110001010010110010110; end
            14'd15448 : begin out <= 64'b0010100010111111001010001110110110101011011111110010100101011011; end
            14'd15449 : begin out <= 64'b1010010010111100101001110000110010100100100011101010101010111011; end
            14'd15450 : begin out <= 64'b1010101011010011001010001000011100101000000001110010101110101001; end
            14'd15451 : begin out <= 64'b0010011100110110001010100111110100101001000111111010011111000011; end
            14'd15452 : begin out <= 64'b0010000001000010001011000000000000101001101111011010100000010110; end
            14'd15453 : begin out <= 64'b1010100010110100001010000100001010011010010011101000011111110000; end
            14'd15454 : begin out <= 64'b1010100111100101101001100000001110101011111000110010101000111011; end
            14'd15455 : begin out <= 64'b1001101000000111001010001111111010101010110010111010010100100111; end
            14'd15456 : begin out <= 64'b1010001100100010101010010101010100100110111100001010011100101111; end
            14'd15457 : begin out <= 64'b0010100000101111101010111100110110100110111010100010101100000011; end
            14'd15458 : begin out <= 64'b0010100010001100101001110100011110101001001100001010010001100001; end
            14'd15459 : begin out <= 64'b1001101011010010101001001100010100101001101110001010101100010010; end
            14'd15460 : begin out <= 64'b1010010000100110001010101000111110101001011111011010001000110111; end
            14'd15461 : begin out <= 64'b0001110010110101001001101000000110100101101010111010100101011101; end
            14'd15462 : begin out <= 64'b1010010011100110100000000010010000101010000011011010110000001010; end
            14'd15463 : begin out <= 64'b1010100101000011101000111001001010101001111000000010010110111001; end
            14'd15464 : begin out <= 64'b0010001100111110101010100110110100011100001111101010100110110000; end
            14'd15465 : begin out <= 64'b1010101111010111001010101001000000100100000110001001010100101110; end
            14'd15466 : begin out <= 64'b0010011100001111101010101111101010011000011111100010100111111110; end
            14'd15467 : begin out <= 64'b0010101011100011101001111011010000100000111010100010101100011111; end
            14'd15468 : begin out <= 64'b0001110001110100101010101011010110101010001011000010011110110110; end
            14'd15469 : begin out <= 64'b0010100111101111101001000011110100101010111011001010100000100000; end
            14'd15470 : begin out <= 64'b0010000011000101001010011001100110101000100111000010101011001000; end
            14'd15471 : begin out <= 64'b0001111001000110101010110011010000101010100000111010101010100110; end
            14'd15472 : begin out <= 64'b0010101110001110000011101000010000101000011011010010000010111110; end
            14'd15473 : begin out <= 64'b0010101000101100000010011001111110101000001100100010100110100100; end
            14'd15474 : begin out <= 64'b1001110101011101001001110010000100100000001010001001110010111010; end
            14'd15475 : begin out <= 64'b0010001111011110001010101001010010100101000000001010101101101110; end
            14'd15476 : begin out <= 64'b0010100110110011001010101010111110011111110011011010101010111110; end
            14'd15477 : begin out <= 64'b0010001000011101101001011000100100100100110101010010011011101011; end
            14'd15478 : begin out <= 64'b1001100001011011001001100000111100100001111111000010100100001001; end
            14'd15479 : begin out <= 64'b1010101101101100101010101001000010100101111101010010011011011011; end
            14'd15480 : begin out <= 64'b1001000100110111001000010000001100101001010000100010101011010111; end
            14'd15481 : begin out <= 64'b0000111011110111101010101010010110101011001010101010100101111000; end
            14'd15482 : begin out <= 64'b1010100000111111100111111110101100101000001101010010101001110011; end
            14'd15483 : begin out <= 64'b1010011111001010101010110000010010101001100100100010011100110000; end
            14'd15484 : begin out <= 64'b0010101000011011101000110001111100101000111101100010100011110001; end
            14'd15485 : begin out <= 64'b0010101101100000101010100000111010100001001100101010100101001101; end
            14'd15486 : begin out <= 64'b0001000100001010101010011101010000101000011100001010010011111000; end
            14'd15487 : begin out <= 64'b1000110110001110001001111001011010100100110100110001101101010101; end
            14'd15488 : begin out <= 64'b0010101110010001101001110111000110101000110011010010101010010001; end
            14'd15489 : begin out <= 64'b1010011110110011001001101101110110011101000000001010100101110100; end
            14'd15490 : begin out <= 64'b1010010000001111000100101100100000100101100001110010011001111110; end
            14'd15491 : begin out <= 64'b1010010011010011101010001111011010100010101101010010100100010111; end
            14'd15492 : begin out <= 64'b1010011010001011001010000000100000101010010101111010000011110000; end
            14'd15493 : begin out <= 64'b1010100101010101000101011011101100101001001111001010011010110010; end
            14'd15494 : begin out <= 64'b0010001000011111101001110011100000100110110111101010011111011111; end
            14'd15495 : begin out <= 64'b0010011101110010101010110010000100101000010111000010001010011011; end
            14'd15496 : begin out <= 64'b1010000110110111101010101110011010100011111000001001101111100001; end
            14'd15497 : begin out <= 64'b0010000000111111101010100110111100100111110111001010100011011111; end
            14'd15498 : begin out <= 64'b0010011000101010001001010110011110101010110001111010000011100000; end
            14'd15499 : begin out <= 64'b1010100100101010001001001101100110011111001100011010100000001000; end
            14'd15500 : begin out <= 64'b0001110101001001101001110001110110100010110100100010011111111001; end
            14'd15501 : begin out <= 64'b1010011010110000001001100010110110101010010001100010100111101110; end
            14'd15502 : begin out <= 64'b1010101100000001100111101011011100101001101110011010011000100011; end
            14'd15503 : begin out <= 64'b1010101110001110001010101111100010010100100100011010100011011011; end
            14'd15504 : begin out <= 64'b1010101110000011001001101001000010100101011010110010010011001110; end
            14'd15505 : begin out <= 64'b1010100001000100001001101111001010101011010111011010010010010111; end
            14'd15506 : begin out <= 64'b1000110101010010101000100111100000100011110010000010101100000010; end
            14'd15507 : begin out <= 64'b1010100101110001101011000000110010100101101000110010101010110011; end
            14'd15508 : begin out <= 64'b1010100110011000001010011011111010101011010111000010101011101001; end
            14'd15509 : begin out <= 64'b1010100110100101001001101110110100101010010010011010101111001011; end
            14'd15510 : begin out <= 64'b0010101000000000001010100111001000100101100011011010010010001110; end
            14'd15511 : begin out <= 64'b1010101101000111000110011110000000101010000111111010101110101110; end
            14'd15512 : begin out <= 64'b1010010011000101101001011111001000011000001100110010101110100100; end
            14'd15513 : begin out <= 64'b1010001100000001001010101010100110100100000101001010010000111010; end
            14'd15514 : begin out <= 64'b1010011011111000101010100110110010101001110101011010101010100100; end
            14'd15515 : begin out <= 64'b1010101100011110101010101111100100100010110110111010101101101010; end
            14'd15516 : begin out <= 64'b1010101111011011101000100111111100100110111000111010011110111100; end
            14'd15517 : begin out <= 64'b1010100111100110001001110111011100011110000101110010100101111110; end
            14'd15518 : begin out <= 64'b0010100101010010101010011010100110101000110100000010101110011110; end
            14'd15519 : begin out <= 64'b0010000110111000101010001000001100100101111101110010101001100111; end
            14'd15520 : begin out <= 64'b0010101011010111001010010101010110101001111001001010100010001101; end
            14'd15521 : begin out <= 64'b1010100010101111001000100000111100100100101110010010011101110010; end
            14'd15522 : begin out <= 64'b0001110110110001001010110000011000011101101011011010101001111100; end
            14'd15523 : begin out <= 64'b0001110100001101101010100110010110100111010110110010110000000011; end
            14'd15524 : begin out <= 64'b0010101011000110101000010000010110100000100010011010101110110101; end
            14'd15525 : begin out <= 64'b0010010110010100001010000101101100100000110101000001001000001100; end
            14'd15526 : begin out <= 64'b0010010110111101101010100010000000101010100000010010101111110101; end
            14'd15527 : begin out <= 64'b1010011100000001001010000000111110100001000110011010001000011101; end
            14'd15528 : begin out <= 64'b1010011000110100001010101001110000101011011001101010101011011100; end
            14'd15529 : begin out <= 64'b0010100000101110101000110111001100011110010001000010101100100100; end
            14'd15530 : begin out <= 64'b1010100100100001101001001011011000010110111000001010101000110000; end
            14'd15531 : begin out <= 64'b1010101001010100001000100110010110100010101110110010101011000001; end
            14'd15532 : begin out <= 64'b1010010111110101000101111000111010010100001000110010100011111101; end
            14'd15533 : begin out <= 64'b0010011101110111101001100111001000101000011110000010101001111001; end
            14'd15534 : begin out <= 64'b0010000011110010101010010101001000101100000001000010011001010100; end
            14'd15535 : begin out <= 64'b1010101111000111000101110000011010101010110110111010001000100101; end
            14'd15536 : begin out <= 64'b0010010110010101000111011100110000010101000011100010100010100001; end
            14'd15537 : begin out <= 64'b1010101000010111001010000100010000101000111001100010101111100011; end
            14'd15538 : begin out <= 64'b0010010111110010001010100100011010101010110101011010000010101111; end
            14'd15539 : begin out <= 64'b1010101011000000001010001010010010011110000111010010011010011111; end
            14'd15540 : begin out <= 64'b0001110101101001101001111100101110101011001010110010100001000110; end
            14'd15541 : begin out <= 64'b1010100110001011001000001011011000100110010000100010100000010101; end
            14'd15542 : begin out <= 64'b0010010001001011101000011111011010101011011011010010010000110100; end
            14'd15543 : begin out <= 64'b0010101110011001101000001000111100101011001011101010000000101001; end
            14'd15544 : begin out <= 64'b1001111011110110001010001101100010011110001000010010010010101011; end
            14'd15545 : begin out <= 64'b1010101101000111001001101111100010101000000001101010100000011110; end
            14'd15546 : begin out <= 64'b0010100111010010001000011001101000101000000100111010000101011100; end
            14'd15547 : begin out <= 64'b0010010111101001001010101010011010101010100110000010100011011000; end
            14'd15548 : begin out <= 64'b0010001100000110101001011001111100101001110001111010011100001111; end
            14'd15549 : begin out <= 64'b1010101011100010101001111001011010101011010100000010100001100110; end
            14'd15550 : begin out <= 64'b1010010111011000101010011111101110100011111100000010000111001011; end
            14'd15551 : begin out <= 64'b1010100100011010001010001111110010011111000011101010101111001100; end
            14'd15552 : begin out <= 64'b1010100100010000001011000010110100101000000011011010101110000001; end
            14'd15553 : begin out <= 64'b0010101001011001001010100000111010101001001000010010101110001000; end
            14'd15554 : begin out <= 64'b0010101111111010101010010010010110101010101111111010101101000100; end
            14'd15555 : begin out <= 64'b0010001101001101001010111111100100011101000010111010101011011111; end
            14'd15556 : begin out <= 64'b1010011101101011101000100101101110100101001001010010000001101101; end
            14'd15557 : begin out <= 64'b1010001010011111101001110100101000100101010000100010001111100110; end
            14'd15558 : begin out <= 64'b1010010010001000101001101000111010100000100011111010101111101000; end
            14'd15559 : begin out <= 64'b1010101100011100000101110101100100101010011101110001110100100101; end
            14'd15560 : begin out <= 64'b0010011111000101101010010111010100100000011111110010101111011010; end
            14'd15561 : begin out <= 64'b1010100100100110100101010001110000101011000010110010101100101010; end
            14'd15562 : begin out <= 64'b0010101101000100000111111101011010101011110010100010001010000100; end
            14'd15563 : begin out <= 64'b1010100110010100001001111100010100101001111111101010101010100011; end
            14'd15564 : begin out <= 64'b0001101110100111001010000100101100100010111000011010101001101110; end
            14'd15565 : begin out <= 64'b1010101011100010101001111110001100001100010011000010100010101100; end
            14'd15566 : begin out <= 64'b0010101011001111101001101001100110101011110100010001111010111101; end
            14'd15567 : begin out <= 64'b0001110101001011101001001011011010101010110000100010100000011010; end
            14'd15568 : begin out <= 64'b1010100010010111101010101001011100100111101111000010000110111111; end
            14'd15569 : begin out <= 64'b0010100011011100101000110110111010100101000110011010100101001101; end
            14'd15570 : begin out <= 64'b0010100110100000101010100101100000101011100100110001101011111111; end
            14'd15571 : begin out <= 64'b0010100101101101101000001010001100100001111100010010100111111011; end
            14'd15572 : begin out <= 64'b1000100111001100001001000111101000011100001101111001100000001001; end
            14'd15573 : begin out <= 64'b0010011101000111101000011100001100101000000000001010101100000101; end
            14'd15574 : begin out <= 64'b0010100111110011101010011001000110011100000101001010100110110000; end
            14'd15575 : begin out <= 64'b0010101010101111101001001010001010101011001000101001110000000011; end
            14'd15576 : begin out <= 64'b0010101111001110001010110000100110100011111011011010100011011000; end
            14'd15577 : begin out <= 64'b1010101100100110101010001010000010100110100010101010100010001100; end
            14'd15578 : begin out <= 64'b1010100011101000001001001100011000100111111111111010001100010111; end
            14'd15579 : begin out <= 64'b0010001000000010001001110000110110101001011010010010011011101111; end
            14'd15580 : begin out <= 64'b0010101101111010101001011110100110101011010110100010010000011000; end
            14'd15581 : begin out <= 64'b1010101010101000000110001011110010000111110110111010010100111000; end
            14'd15582 : begin out <= 64'b1010100010110010001001110010111010100100101010110010001100000011; end
            14'd15583 : begin out <= 64'b1010010110100100001000100100000000100001110010011010010110001001; end
            14'd15584 : begin out <= 64'b0010101011000000001001011010111100100111110100010010001011110101; end
            14'd15585 : begin out <= 64'b1010100101101100100111000110101010101001000010001010101110111000; end
            14'd15586 : begin out <= 64'b1010100111100110101001111010110110010100111101111010101010001110; end
            14'd15587 : begin out <= 64'b0010100101110111000111101010110100101010100111010010100110010110; end
            14'd15588 : begin out <= 64'b1010101010010001001010101000001000100101110111011010001100111000; end
            14'd15589 : begin out <= 64'b1010100010111000000110001001100100101001001011010010001100110101; end
            14'd15590 : begin out <= 64'b1010010011011100101000110011111010101001110000111010011111011011; end
            14'd15591 : begin out <= 64'b1010000100110101000110010100001010101010111000100010101110011101; end
            14'd15592 : begin out <= 64'b1010100010001101001010111110011000101010011011110010110000000111; end
            14'd15593 : begin out <= 64'b0010010010010100001001000011111100101011100110010010010111010010; end
            14'd15594 : begin out <= 64'b0010010000100011101010111110001100101001000111011010100101010011; end
            14'd15595 : begin out <= 64'b1010101100011111101000011111001100101010111110110010011111100001; end
            14'd15596 : begin out <= 64'b1010000000000101101000111111000010101001110100101001111101100110; end
            14'd15597 : begin out <= 64'b0010011101101011001001000000001010101011010100100010101010011010; end
            14'd15598 : begin out <= 64'b0010101010100100001000010101100000101000110100001010011101001000; end
            14'd15599 : begin out <= 64'b1010011110011110000110111001101010101000101111111010010010101000; end
            14'd15600 : begin out <= 64'b0010101011001111101010000000000000101010111111111001111100100100; end
            14'd15601 : begin out <= 64'b0010101001001001001010100101000010011100101110100010011001011001; end
            14'd15602 : begin out <= 64'b0010011001101010000110010000010110100101001010100001100000010101; end
            14'd15603 : begin out <= 64'b1010100001010000101010111011101010100001100101011010011100010100; end
            14'd15604 : begin out <= 64'b0010100011111111001010100111010110101011111000010010000000111010; end
            14'd15605 : begin out <= 64'b0010010001111011101010111100010100101100001010101010010111100110; end
            14'd15606 : begin out <= 64'b1010100010110011100111111010111000100110100101110001110011001111; end
            14'd15607 : begin out <= 64'b1010100010101011101000110010000010011011101000010010101110001110; end
            14'd15608 : begin out <= 64'b0010010101000100101010000011000000000100111111011010101111000000; end
            14'd15609 : begin out <= 64'b1010100110000011001010111001010110101001111010100001110110100011; end
            14'd15610 : begin out <= 64'b1010100110101100100111100001001000100111011100101010100101100011; end
            14'd15611 : begin out <= 64'b1010101101111111001001001111010100101001111010011010100110001001; end
            14'd15612 : begin out <= 64'b0010100000111111001010100000010110101100000010010010101001011100; end
            14'd15613 : begin out <= 64'b1010010010100011101010010001110010100111101000101010010011110111; end
            14'd15614 : begin out <= 64'b1001100111011001001010101011011110101100000000101010101001101010; end
            14'd15615 : begin out <= 64'b1010000010010111101010100100001000101010101011010010011011010010; end
            14'd15616 : begin out <= 64'b1010100011001011001010010011111110101001100111111010010000011101; end
            14'd15617 : begin out <= 64'b1010100010111010001010011000011100101011110010011010101110100110; end
            14'd15618 : begin out <= 64'b1010101001110110001010001001101110100100101000001010100011100010; end
            14'd15619 : begin out <= 64'b1010011100010001000001100101001000101010101100010010000000110010; end
            14'd15620 : begin out <= 64'b0010101010101010101001100000011110101011110111000010101000000101; end
            14'd15621 : begin out <= 64'b1010100100011100101001010001011110101011101100100010010010100111; end
            14'd15622 : begin out <= 64'b1010011001011001001010110101001110101011101101101001111100001000; end
            14'd15623 : begin out <= 64'b0010010100110010001010001010000100100010000110111010101010000001; end
            14'd15624 : begin out <= 64'b0010011110101001000111110000001000100111000000110010011011100111; end
            14'd15625 : begin out <= 64'b0010011101101010001010011010100010100100010100000001010101001101; end
            14'd15626 : begin out <= 64'b1010010001100100101010110110101100100101011000011010101100100010; end
            14'd15627 : begin out <= 64'b1010101100010111001010110110100000100101111110011010101110000101; end
            14'd15628 : begin out <= 64'b0010100010000011100111110011101000101000000011110010010010010110; end
            14'd15629 : begin out <= 64'b1010100011100111001001101111001110101011010001100010010111101110; end
            14'd15630 : begin out <= 64'b0001101000010010000111111000110000100110010100101010100010010001; end
            14'd15631 : begin out <= 64'b0010101101100111101010010001111010100000100011011010100010001101; end
            14'd15632 : begin out <= 64'b1010100100000110000011101101000000100100111111001010010001010001; end
            14'd15633 : begin out <= 64'b1010000011010000001001110101111010100111100101001010100011101111; end
            14'd15634 : begin out <= 64'b1010101000100101000111011010001000101001100101010010000101011011; end
            14'd15635 : begin out <= 64'b0010010110000100000100100110111100011010100100111010100100011100; end
            14'd15636 : begin out <= 64'b1010011010011101100110110111101000100110001010100010101110110001; end
            14'd15637 : begin out <= 64'b0010100110110101001010101101110000101000001111101010010100001010; end
            14'd15638 : begin out <= 64'b0010011101011000101010110100111010100101111010100010100001111111; end
            14'd15639 : begin out <= 64'b1010100001100110101001000001111100100111110001001010100001000101; end
            14'd15640 : begin out <= 64'b0010100111011111101001000101101010100111111101110010010001111010; end
            14'd15641 : begin out <= 64'b0010000100000100001010101010101110101001110010100010101111100001; end
            14'd15642 : begin out <= 64'b1010010101110010100110000001101010101010010101011001010011110101; end
            14'd15643 : begin out <= 64'b1010010011000111101010010111110110101000101011010010001010010100; end
            14'd15644 : begin out <= 64'b1010100001111100101000100010111010101011110111101010100010000101; end
            14'd15645 : begin out <= 64'b0001110100110111001001010111000010101000010011010010101100111111; end
            14'd15646 : begin out <= 64'b0010101011111010001010000101001110011001011100010001110000000110; end
            14'd15647 : begin out <= 64'b0010001011100111101010010001011000101010000000110010100100101011; end
            14'd15648 : begin out <= 64'b0010100101100000100111101001011110100001100010101010101111101100; end
            14'd15649 : begin out <= 64'b1010101101001111001000001101000000011111001001001010100110011101; end
            14'd15650 : begin out <= 64'b0010000111011111001001001000110010101001011100111010100101011111; end
            14'd15651 : begin out <= 64'b1010001100011000001010101100110100101000101010110010011110100101; end
            14'd15652 : begin out <= 64'b1010011111001010001010101010100100011000110011011010010011001011; end
            14'd15653 : begin out <= 64'b1010011110000100101010010100110010101010111011100001111001011111; end
            14'd15654 : begin out <= 64'b1010000101001100001010001010111110101011010001111010010111100000; end
            14'd15655 : begin out <= 64'b1001101111000100001010001010111000011111111011001010101011101111; end
            14'd15656 : begin out <= 64'b0010010101010011001010100000111010001110011001110001110010111001; end
            14'd15657 : begin out <= 64'b1010100111100000101010100101000000011101010010101010010011100111; end
            14'd15658 : begin out <= 64'b1010010100001011101010001111110010100010000011111010011011001011; end
            14'd15659 : begin out <= 64'b1010100100001001101010111111111000101001001110000010100101000010; end
            14'd15660 : begin out <= 64'b1001111110110001000100101000001010001111010000011001111111101101; end
            14'd15661 : begin out <= 64'b0010011011110110001010111010010010101010100111111010100110111100; end
            14'd15662 : begin out <= 64'b0010100111010110001010011110000110101000000111011010101100010101; end
            14'd15663 : begin out <= 64'b0010100011000011001010001000011010100000011110110010101100000011; end
            14'd15664 : begin out <= 64'b0010011100100101001000001011011110101000100000110010100010101101; end
            14'd15665 : begin out <= 64'b0010100111100000101010001101011000101000111101110010011000000110; end
            14'd15666 : begin out <= 64'b1010101101000101100110000101011100100110100010100010010100101000; end
            14'd15667 : begin out <= 64'b0001110101001000101010111011011110101100001010001010011110101000; end
            14'd15668 : begin out <= 64'b0010100011110001100111101110111010101100001001110010010110110110; end
            14'd15669 : begin out <= 64'b1000110101111110101010101111001010100011100110010010101110100000; end
            14'd15670 : begin out <= 64'b1010011111010111000111101000010000101001001001100010001000101111; end
            14'd15671 : begin out <= 64'b0010101100101100101001011101000000101001110110001010101101111101; end
            14'd15672 : begin out <= 64'b1010100111100001001010010001000010100110001111110010001000010011; end
            14'd15673 : begin out <= 64'b1010100011111101001000011001011000101011111000010010011010101011; end
            14'd15674 : begin out <= 64'b0010010011100001101010100001001110011111000110001010101110110000; end
            14'd15675 : begin out <= 64'b1010101000100010001000000110100000100101100100100010101010110110; end
            14'd15676 : begin out <= 64'b0010101000001001100110000111111000100110011110111010000011001101; end
            14'd15677 : begin out <= 64'b0010100101000010101001110101111100100110100100010010010010011101; end
            14'd15678 : begin out <= 64'b0001101111010011101001000110001010100010001100101010011111001100; end
            14'd15679 : begin out <= 64'b0010010111100101001001011000011010101000110011100010100101111010; end
            14'd15680 : begin out <= 64'b1010010110000000101010000011001010100010111001111010010110100011; end
            14'd15681 : begin out <= 64'b0010001001110110101001010001110000101010110100111001100110100011; end
            14'd15682 : begin out <= 64'b1001110110010011101000001101101100101010000100111010010011110001; end
            14'd15683 : begin out <= 64'b1010001111001001100101111010101010101001011001101010011110000011; end
            14'd15684 : begin out <= 64'b1010101101010010101000000101011000010101011011100001110111100101; end
            14'd15685 : begin out <= 64'b0010001100111011001000011100110010100001010000101010010100010001; end
            14'd15686 : begin out <= 64'b0010001011111010001010010001010110101000111010101010011000100001; end
            14'd15687 : begin out <= 64'b1010101000111110001001101111100110100110001010010001111000110000; end
            14'd15688 : begin out <= 64'b0010100101100010101010001100101000101011110100010010001100001000; end
            14'd15689 : begin out <= 64'b1010001011001100101010101110010000010100010000101010001111101100; end
            14'd15690 : begin out <= 64'b0001101100110011001010001010111010100001010000101010100011001100; end
            14'd15691 : begin out <= 64'b0010010111101110001000101010101110101000110101111010101100110001; end
            14'd15692 : begin out <= 64'b1010100000001011000110110100010110100110101110111010101000100000; end
            14'd15693 : begin out <= 64'b1010100100010110101000000100100010101010111010100010100011010000; end
            14'd15694 : begin out <= 64'b0010001010110101101000010011011000101000101000101010101011000100; end
            14'd15695 : begin out <= 64'b0010101010010111100111011101110000101011100101101010100110000111; end
            14'd15696 : begin out <= 64'b0010100110010010001000100100001010101100000100111010011010100011; end
            14'd15697 : begin out <= 64'b0010101000010000101010101000111000011110110001101001110011100001; end
            14'd15698 : begin out <= 64'b1001011010011011001010010010100010101010011111100010010000100100; end
            14'd15699 : begin out <= 64'b1001101000001111101010000010001000101000010001111010010111111110; end
            14'd15700 : begin out <= 64'b0010000001001000101010001001000110100111100110011010011101010001; end
            14'd15701 : begin out <= 64'b1010011000110111101010001111010010010111101111100001111100000000; end
            14'd15702 : begin out <= 64'b0010011000111101001010010011010010011111111001010010100000110110; end
            14'd15703 : begin out <= 64'b0010010001111110001000000000000100100111100000110010011001101011; end
            14'd15704 : begin out <= 64'b0010100101101000001010100100001110101000111101011001101101000010; end
            14'd15705 : begin out <= 64'b0010000101100101101010100111101000101011100001011010101001111010; end
            14'd15706 : begin out <= 64'b0010100100000001101010110111010010000111100100111010011000100101; end
            14'd15707 : begin out <= 64'b1010010010111000001010001110101100100110010010111001111101101010; end
            14'd15708 : begin out <= 64'b0010000110001000001010110001001000101010000000000001101100100101; end
            14'd15709 : begin out <= 64'b1010100011110000001010001111000000101010111110010010101111010111; end
            14'd15710 : begin out <= 64'b1010000111101111101000111001100000101010110101101010010100111000; end
            14'd15711 : begin out <= 64'b0010100000101110001001100100101100101000010000110010001001101000; end
            14'd15712 : begin out <= 64'b1001110000011111001001010111000010101011110111011010100001101001; end
            14'd15713 : begin out <= 64'b1001110000110100001001111001011000100101001011101010010100110001; end
            14'd15714 : begin out <= 64'b1001001001000000101010111111100000100111101010101010011001011101; end
            14'd15715 : begin out <= 64'b1010000100111010000110000001110000101011001111010010101011100110; end
            14'd15716 : begin out <= 64'b1010001111001101101010001111111100100010001110010010010110111010; end
            14'd15717 : begin out <= 64'b0010101010010111001000001001101100100010110000110010101100110111; end
            14'd15718 : begin out <= 64'b1010100001100000001010101001100000100000100010100010100011101000; end
            14'd15719 : begin out <= 64'b1010011110110000101010000110000000101001011001000010100000010001; end
            14'd15720 : begin out <= 64'b1010011010001010001010010000010100101010010011111010101110011100; end
            14'd15721 : begin out <= 64'b0010101000100010001010001001001110100111000101001010101101110111; end
            14'd15722 : begin out <= 64'b1001101010100001001001110101101000101011010111011010100100000011; end
            14'd15723 : begin out <= 64'b1001010111110110000110011111111010101011010010001010101100010111; end
            14'd15724 : begin out <= 64'b1010100111100011101010111001010000100000010101111010100010110000; end
            14'd15725 : begin out <= 64'b0010100001011001101000110101010010101011001001100010100011011110; end
            14'd15726 : begin out <= 64'b0010100000111011100111010010011100100000011000111010100110000010; end
            14'd15727 : begin out <= 64'b1010001011010101101010001101100110100110100100010010100110010011; end
            14'd15728 : begin out <= 64'b1010101010001011101001101010100000101000010101110001101000011101; end
            14'd15729 : begin out <= 64'b1010101000010000101010010000100100011110010001001010100100100001; end
            14'd15730 : begin out <= 64'b0010101010001010101010101000101010010110100001101010100111111110; end
            14'd15731 : begin out <= 64'b1010000000010011001001001100010010100101101110110010100100011011; end
            14'd15732 : begin out <= 64'b0001011101001001001010100000101110011100101101100010100110101100; end
            14'd15733 : begin out <= 64'b1010101010010100001001001101100100101000101110001010000011001011; end
            14'd15734 : begin out <= 64'b0010010111100110101010001101001110100101011101000010100011101100; end
            14'd15735 : begin out <= 64'b0010100100101110001000110100100010100011101001111010001011101000; end
            14'd15736 : begin out <= 64'b1010011100100001101010001111000010100001000010101010101101110100; end
            14'd15737 : begin out <= 64'b1010010101010101001001101011000100101010000000110001101111111000; end
            14'd15738 : begin out <= 64'b0010101001000010101000000100110010101001010110100010010110101000; end
            14'd15739 : begin out <= 64'b1010101100110000001001110101010100100110111001000010101110000001; end
            14'd15740 : begin out <= 64'b0000001000011110101010100000111110100011010100111010100010001110; end
            14'd15741 : begin out <= 64'b1010001101000110100111010011000000100000110101101010010111110001; end
            14'd15742 : begin out <= 64'b0010010111000001101010101011110010101000011100111010011110011101; end
            14'd15743 : begin out <= 64'b0010101100010000101000101001110110100010100100100010010100000111; end
            14'd15744 : begin out <= 64'b0010001101110101101010100010000100010111101100010010100101011011; end
            14'd15745 : begin out <= 64'b0001110011101011001001000011010000100111001100000010101010010000; end
            14'd15746 : begin out <= 64'b1010100011001011101010000101011110100111010101100010011000011001; end
            14'd15747 : begin out <= 64'b1010000101000110101010101100001100101010000101100010000111000001; end
            14'd15748 : begin out <= 64'b0010101110110101101010100011011110100101001010100010010101001010; end
            14'd15749 : begin out <= 64'b0010100000011001100111010010000100100111001010001010010110110000; end
            14'd15750 : begin out <= 64'b1010000101010011101010101000011100100000110000010010001010011010; end
            14'd15751 : begin out <= 64'b1001110100000111101001000001010010011110101011011010011100001101; end
            14'd15752 : begin out <= 64'b0010101000000100101000110110011110101000010101111010101001011111; end
            14'd15753 : begin out <= 64'b0010101000011110101000101001101000100101101001000010011001110001; end
            14'd15754 : begin out <= 64'b1010101010100100001001100110011000101011011101010010101111010000; end
            14'd15755 : begin out <= 64'b0010100110111011001000100010011010100101100000001010100101110100; end
            14'd15756 : begin out <= 64'b1010010100110001101001011101001010100111110010011010001001101110; end
            14'd15757 : begin out <= 64'b0001111110100001001000001011001110101011101001111010001010101001; end
            14'd15758 : begin out <= 64'b0001000001110111100111100111110110100111111001111010100001011010; end
            14'd15759 : begin out <= 64'b1010001111011110101010100100011110101011011111111010100100100011; end
            14'd15760 : begin out <= 64'b0010010001100110001010000000101100100111111111110010001000111110; end
            14'd15761 : begin out <= 64'b0010100010000000001001011101010100101001111011001010100100010010; end
            14'd15762 : begin out <= 64'b1010101010011001101000110011001000100100010000110010101110110001; end
            14'd15763 : begin out <= 64'b1010100000011100001001101000111110100010011011111010100100001010; end
            14'd15764 : begin out <= 64'b0001101100010010101001101000011000101001100100101010100100010111; end
            14'd15765 : begin out <= 64'b0010100011110111001010010001111000100011101000110010000101111000; end
            14'd15766 : begin out <= 64'b1001101111010101101010011101110100100101100011101010101101100010; end
            14'd15767 : begin out <= 64'b0001111101001010001001001111111110100010000000000010011010001110; end
            14'd15768 : begin out <= 64'b0010101011000001001010100001111110101001000010101010001000000000; end
            14'd15769 : begin out <= 64'b0010100011110110001001100110101000100010011100100010101000011101; end
            14'd15770 : begin out <= 64'b0010100011100010101010100010111000101011000001001010010001001101; end
            14'd15771 : begin out <= 64'b1010101001101001101010011110001110101010110101101010100000101110; end
            14'd15772 : begin out <= 64'b0010001100001010001010100110101010101001011000000010101101000000; end
            14'd15773 : begin out <= 64'b1001110100100111101000110100110110100100110001111010001100100111; end
            14'd15774 : begin out <= 64'b1010101001010011001010011011001010101001111001001010100100010000; end
            14'd15775 : begin out <= 64'b0010010001100101001000001010011100101011100111000010010111111100; end
            14'd15776 : begin out <= 64'b1010101101110111101001100110010110101011101001001010100010001110; end
            14'd15777 : begin out <= 64'b1010100010111011100111101101011000100100010110001010010010001001; end
            14'd15778 : begin out <= 64'b1010010110011000100111011011100100101000111011101010100000010010; end
            14'd15779 : begin out <= 64'b1010100010010000101010100011010000101001000011001010101101111010; end
            14'd15780 : begin out <= 64'b1010000110010101001010101101010010011110101101010010010100001110; end
            14'd15781 : begin out <= 64'b0010101110101110001010000001111000100101110011111010001111100101; end
            14'd15782 : begin out <= 64'b0001100111010111101010111101000100101001100011101001100001011100; end
            14'd15783 : begin out <= 64'b1010010100001100001001000011110100100100001011010010100110111111; end
            14'd15784 : begin out <= 64'b0001000110001111001010010101011010011010111101101010011010110000; end
            14'd15785 : begin out <= 64'b0010011011100010101010101101001010101011101111000010100001111100; end
            14'd15786 : begin out <= 64'b1010000001011111001010010100110100101010001111100010101111011011; end
            14'd15787 : begin out <= 64'b0010011011011110101010010011111010101000000000010010100000110000; end
            14'd15788 : begin out <= 64'b1010101111011000001010101100100000101010001101110010100111110010; end
            14'd15789 : begin out <= 64'b1010100111011100001010100110100110101001101111101010100110000111; end
            14'd15790 : begin out <= 64'b1010100010100000001010000001110110100110110100000010011000110000; end
            14'd15791 : begin out <= 64'b0001010110010110001010011000111010101010001101000001101111000101; end
            14'd15792 : begin out <= 64'b1010101100010100001001111101101100101000000010001010011101010110; end
            14'd15793 : begin out <= 64'b0010100000100010101001001101011100101011010111101010101111111011; end
            14'd15794 : begin out <= 64'b1010101011001110001010001000111010100111010111111010101111000010; end
            14'd15795 : begin out <= 64'b0010101010110011001010011011010010101000111101110010100010011110; end
            14'd15796 : begin out <= 64'b1010001010010110001010010010111110100100100011101010011010010111; end
            14'd15797 : begin out <= 64'b0010001010111100101010101011111000100111100100110010000011101010; end
            14'd15798 : begin out <= 64'b0001111111011110101010101001001000101000100101101010101001000001; end
            14'd15799 : begin out <= 64'b0001110100011011001010000010010000101001110010011010010111101101; end
            14'd15800 : begin out <= 64'b0010101111100110001010111001100100100111100011010010011010111010; end
            14'd15801 : begin out <= 64'b1010101110001110001010111011011000100101011010000010100000101101; end
            14'd15802 : begin out <= 64'b0010100110011101101010001010100110101001101000001010101000001100; end
            14'd15803 : begin out <= 64'b0010001011111101001010101010010100101000010000010001100000110010; end
            14'd15804 : begin out <= 64'b0010101111111110101001000000011100011011011001000010001000110001; end
            14'd15805 : begin out <= 64'b1001111101101000000111010110110000101010000011101010010010101010; end
            14'd15806 : begin out <= 64'b1010101100110110101000010011110100101000001000100001111000111101; end
            14'd15807 : begin out <= 64'b1010101010100000001001110111100010101010100111011010100101000110; end
            14'd15808 : begin out <= 64'b1010101000001110001010110101101010101011011001110010101011100101; end
            14'd15809 : begin out <= 64'b1010011110110111101010011010111100101011001000000001110111101110; end
            14'd15810 : begin out <= 64'b1001110101111011001010101100001110100101001111000010100011010110; end
            14'd15811 : begin out <= 64'b1010000111001101001001101000000110010000100001001010100011101101; end
            14'd15812 : begin out <= 64'b0010101000100100001001011100111010101011000000110010100000011110; end
            14'd15813 : begin out <= 64'b1010100001100110101010101101110010011101111100100010101110000101; end
            14'd15814 : begin out <= 64'b1010011111111011101010110011111110100110010001100010100001010100; end
            14'd15815 : begin out <= 64'b0010010110010001001000101010111010101001011111010010101110111010; end
            14'd15816 : begin out <= 64'b1010101011011000101000111110111110100111100100010010101001011111; end
            14'd15817 : begin out <= 64'b1010101111000110000111110000100010100010010100100010101011100011; end
            14'd15818 : begin out <= 64'b1010100100101111001010011111011000100111010101101010011001001001; end
            14'd15819 : begin out <= 64'b1010101101101001001010000000011010100111010111100010101101011110; end
            14'd15820 : begin out <= 64'b1001100001111011101010111011000100101011101101000010100000011010; end
            14'd15821 : begin out <= 64'b1010101101010010101001001000101110100111111000001010100101110001; end
            14'd15822 : begin out <= 64'b0001101010000011001000011110001110001000011100000010010110000010; end
            14'd15823 : begin out <= 64'b0010001010000111100111011000111100101000011000010010101110011010; end
            14'd15824 : begin out <= 64'b1010011101011111101000100010010000011001001100000010101011101111; end
            14'd15825 : begin out <= 64'b0001110100001010001010101001010000101001000011011010010100000100; end
            14'd15826 : begin out <= 64'b0010100100110100001001101000010100100001001011101010011100011100; end
            14'd15827 : begin out <= 64'b1010101101111100101010010001101000100101101110101010101101100000; end
            14'd15828 : begin out <= 64'b1010101010011010001010010100011000011100110010010001110111100100; end
            14'd15829 : begin out <= 64'b1010100010010111001001101101010110101010101111101010100010111100; end
            14'd15830 : begin out <= 64'b1010101110110001101001111010101010100110101101110010101010011011; end
            14'd15831 : begin out <= 64'b1010011110100000101010011010000100101001110110011010100110001001; end
            14'd15832 : begin out <= 64'b1010011010110011001010111110111110100110100000101010100000000101; end
            14'd15833 : begin out <= 64'b0010000110011100001001110101111000100000011111011010101001101001; end
            14'd15834 : begin out <= 64'b0010100110111000001001001110011000101010010101011010010000000100; end
            14'd15835 : begin out <= 64'b1010000000111100100101111110000000101000100111110001110101010111; end
            14'd15836 : begin out <= 64'b0010100010111001001010010010100000100110001000001010100011001110; end
            14'd15837 : begin out <= 64'b1010011110000110101001011111000010011011000000011010101111011010; end
            14'd15838 : begin out <= 64'b1010001011101011001001110011010000101001001000100010101000000011; end
            14'd15839 : begin out <= 64'b0010011010011110101010101100101100101000010011010010100101110110; end
            14'd15840 : begin out <= 64'b1010000111000110001001000101001100100001101111000010100011101111; end
            14'd15841 : begin out <= 64'b0010010010101000101010010100101100100101110111010010101011110010; end
            14'd15842 : begin out <= 64'b1010101011011010001010110101101010101011100100010010101010101001; end
            14'd15843 : begin out <= 64'b0010011010011100001010100010000110100101111001010001011010000101; end
            14'd15844 : begin out <= 64'b0010000011000111101000101001011000100111010010111010101100000101; end
            14'd15845 : begin out <= 64'b1010101111001001101001010110001100101001100001101001101001101000; end
            14'd15846 : begin out <= 64'b1010100110011111101010100101001010101011100110001010001010011111; end
            14'd15847 : begin out <= 64'b0010101111011110101010100001111010100001111100000010010000001111; end
            14'd15848 : begin out <= 64'b0010101010100111101000000110010010100111110111100010001000001110; end
            14'd15849 : begin out <= 64'b0010011000110110001010101001110000101000000111100010010000001001; end
            14'd15850 : begin out <= 64'b0010101110100000101000011011101010101001110111101010001001101101; end
            14'd15851 : begin out <= 64'b0001111110001100101001110011111010100110001011001010000001111110; end
            14'd15852 : begin out <= 64'b0010000001101111101001101101000110101011100011011010100010010110; end
            14'd15853 : begin out <= 64'b1010101011101101101010101010110100101010000101000010100001010010; end
            14'd15854 : begin out <= 64'b1001010010000111100101010010001100101001010111100010011101111001; end
            14'd15855 : begin out <= 64'b1001110011110010101010111011000000100110101000111010010110000011; end
            14'd15856 : begin out <= 64'b1010101001101100001010010100000110101100001001101010100011110100; end
            14'd15857 : begin out <= 64'b1001111101001010001000111110101000100011111111100010100100010000; end
            14'd15858 : begin out <= 64'b0010101011110111001001000101001110101001011101010010100001000000; end
            14'd15859 : begin out <= 64'b1010011000010100101010011111111000001101110011100010100110001110; end
            14'd15860 : begin out <= 64'b0001101000001010000110010100001110100111000100111001011010110111; end
            14'd15861 : begin out <= 64'b1010011111100101001001111111110000101001001100001010100010011100; end
            14'd15862 : begin out <= 64'b1001110000000011001001000011111100101001000011111010010101011000; end
            14'd15863 : begin out <= 64'b1010101001111001000110011001001000100110000000000010100011010100; end
            14'd15864 : begin out <= 64'b0010100110101110101001001011010110101011110100010010000000011000; end
            14'd15865 : begin out <= 64'b1001010100100011001001000101100000101011001110101010010101110100; end
            14'd15866 : begin out <= 64'b0010100110100101101001111011101110101010111010011010101110110111; end
            14'd15867 : begin out <= 64'b0010101001111100101001001110001100100101100101010010101111110111; end
            14'd15868 : begin out <= 64'b0010100101100000001010011100100110100010111110100001111110001011; end
            14'd15869 : begin out <= 64'b1010010010101000001000110111111100100100110101000010011110111001; end
            14'd15870 : begin out <= 64'b0010001000100101001001111110101010101000100100100010100111110010; end
            14'd15871 : begin out <= 64'b1010001110111111001010010100011100100110011001010010100011110001; end
            14'd15872 : begin out <= 64'b0010101001001001101010011101010100100110001010101010100100010101; end
            14'd15873 : begin out <= 64'b0010100011110111100110101111101010101001000100111010101100110001; end
            14'd15874 : begin out <= 64'b0010101000010000001000110101000010101010110011111010010000100000; end
            14'd15875 : begin out <= 64'b1010100110111100101000001001101100101001010001100010110000001011; end
            14'd15876 : begin out <= 64'b0010100100011010101000111010100110011100101011001010011101101100; end
            14'd15877 : begin out <= 64'b1010101001100111001001100100110000101001000100001010100011101001; end
            14'd15878 : begin out <= 64'b0010100010010100101010001000010100100101111001101001100110010011; end
            14'd15879 : begin out <= 64'b1010101011010000101001110000101010101000110001001010000011001001; end
            14'd15880 : begin out <= 64'b1010100011100100101010110001101110101001001100111010011101001110; end
            14'd15881 : begin out <= 64'b0010100101111001101011000000011100101000001011110010100010011011; end
            14'd15882 : begin out <= 64'b0010011011111110101010110000101010010000010111101010100110111000; end
            14'd15883 : begin out <= 64'b1010101010011110101010011100100010101010100010110001110111100011; end
            14'd15884 : begin out <= 64'b1010010111010101000111001100100000100100111111110010101000110111; end
            14'd15885 : begin out <= 64'b1010101101011000101010000110101100101010111010011001111101000111; end
            14'd15886 : begin out <= 64'b0010101000100000000111100001110010100001100110111010010110101110; end
            14'd15887 : begin out <= 64'b1010001011010101101000100100111010101000101100011010100111011011; end
            14'd15888 : begin out <= 64'b1010010001011001001001011000110100101010111100011010011110011001; end
            14'd15889 : begin out <= 64'b1010100110000110001001011011000100011100101000101010000111101001; end
            14'd15890 : begin out <= 64'b1010000100110010001010010010010010101001001010101010101011000100; end
            14'd15891 : begin out <= 64'b0010100010010101001010010010010000100011001010000010010001101000; end
            14'd15892 : begin out <= 64'b1010011111101111001000110000101100101000111101010010100010000111; end
            14'd15893 : begin out <= 64'b0010101011110101001010111111001100101000011011010010100100101011; end
            14'd15894 : begin out <= 64'b0010010011011010101010111100001010101010001000001001000010000011; end
            14'd15895 : begin out <= 64'b0010101011010011101001100011000110100100010000010010010111001110; end
            14'd15896 : begin out <= 64'b1010100111100110101001011001110010101010101011011010100010110001; end
            14'd15897 : begin out <= 64'b0001111100110011101010010100110110011110001011111010101010100011; end
            14'd15898 : begin out <= 64'b0010100011011010001010111001110010100101111001001010101001100100; end
            14'd15899 : begin out <= 64'b1010010001101011101010101100101110101001011000100010100011110100; end
            14'd15900 : begin out <= 64'b1010101010000010001010000110000010100100110100100010101000110000; end
            14'd15901 : begin out <= 64'b0010011101100101101001111110110000010111010111010010000011000001; end
            14'd15902 : begin out <= 64'b0010101110110011101010010000010100100110010101101010100111000001; end
            14'd15903 : begin out <= 64'b0010100001010001001010011001010000101001110101010010000101101011; end
            14'd15904 : begin out <= 64'b1010011010001111101001111101111100100100110010110010010000110101; end
            14'd15905 : begin out <= 64'b1010000110001101101010011000101110101001111001001010010100110110; end
            14'd15906 : begin out <= 64'b1001110011000011101010010001011010100111001000100010011111111111; end
            14'd15907 : begin out <= 64'b0010001010111110101010010110101100101011100001111010011100011011; end
            14'd15908 : begin out <= 64'b1010100010101110001010001110010110101000100101110010101001011001; end
            14'd15909 : begin out <= 64'b1010100111011001001010111100100100101010111101100010101010011101; end
            14'd15910 : begin out <= 64'b0001011100100100001010011000011000100111101110101010101111111100; end
            14'd15911 : begin out <= 64'b1010010010010010101001000101010010100101101000010001111000110101; end
            14'd15912 : begin out <= 64'b0010011000010001001001111000110000010100110011111010100100110101; end
            14'd15913 : begin out <= 64'b1010100111101111101010001011011100100100110001000010011011111011; end
            14'd15914 : begin out <= 64'b1010011110010100001001111101101010100111100100111001110100000111; end
            14'd15915 : begin out <= 64'b0010101001010110001010101100111010101011001010011010110001000100; end
            14'd15916 : begin out <= 64'b1010010110001010001001000100110010101010110101100010101111111010; end
            14'd15917 : begin out <= 64'b0010100001110000101010011001000000101010011100011010011000111110; end
            14'd15918 : begin out <= 64'b0010000001100111101010000011100010011101100001111010011011010000; end
            14'd15919 : begin out <= 64'b1010010011010001100111011010101010100101000001010010101111001111; end
            14'd15920 : begin out <= 64'b0010101011000111001000001100111000011110100110111001101101111110; end
            14'd15921 : begin out <= 64'b1010101001110110001000100000100010100101011101001010100010111001; end
            14'd15922 : begin out <= 64'b1010101010101111001010110001001100100011101100110010101100001111; end
            14'd15923 : begin out <= 64'b1010101101101101101010001011101110101000001001000010001111111001; end
            14'd15924 : begin out <= 64'b1010101100100011001010110111100110011100011110001010011111011101; end
            14'd15925 : begin out <= 64'b1010010010110010001001101010100100101010101001001000101110101110; end
            14'd15926 : begin out <= 64'b1010100100010011001010000010000100101001110000101010010001010011; end
            14'd15927 : begin out <= 64'b0001011100010000101011000000001110011110111110110010011001101011; end
            14'd15928 : begin out <= 64'b1010010111010101101001011100100100101010111000101010010010110101; end
            14'd15929 : begin out <= 64'b1010010111111111101010100110000010100111101000111010011010001010; end
            14'd15930 : begin out <= 64'b0010101011111100001010100110100100100011011001010010010100001110; end
            14'd15931 : begin out <= 64'b0010100001110101101010000101010110101000011100010010101110100010; end
            14'd15932 : begin out <= 64'b1010000111010000001000011011111100011111010011101010100001111100; end
            14'd15933 : begin out <= 64'b0010011101010011101000111111111110100101000001110010100100011110; end
            14'd15934 : begin out <= 64'b0010011001001110101010100001100100101000100101001010100110101100; end
            14'd15935 : begin out <= 64'b0010011001100101001001111111111110100000000111010010101110010010; end
            14'd15936 : begin out <= 64'b0010010100111010101001011110110100101001001100111010101001101100; end
            14'd15937 : begin out <= 64'b1010001010001001101000100111111100100100101100100010100101100010; end
            14'd15938 : begin out <= 64'b1010010110101110001010100011100110011010000001111010101011110110; end
            14'd15939 : begin out <= 64'b1010101100110011101001100100101110100100110111110010100101010100; end
            14'd15940 : begin out <= 64'b1010000010000110101001011110110100101011110110001010011110101101; end
            14'd15941 : begin out <= 64'b1010100101100011001010011101110100011010010011111010101111110000; end
            14'd15942 : begin out <= 64'b1010101100001100101000011101100010011101111100000010100000010001; end
            14'd15943 : begin out <= 64'b0010001100010001101000011111011110101001101011011010100011001011; end
            14'd15944 : begin out <= 64'b0010001011001100101010010110001100101001101100110010100011000101; end
            14'd15945 : begin out <= 64'b1000000111101100101001011010101100101000010011101010101011111010; end
            14'd15946 : begin out <= 64'b1010010000110111001000111101111100101000011011000010100011001001; end
            14'd15947 : begin out <= 64'b1010001001110101100111101111100100100000001101001010101000100001; end
            14'd15948 : begin out <= 64'b0010011001100001101010001000101010101011100011000001011101110000; end
            14'd15949 : begin out <= 64'b1010001100011111101010100101101110010100001100000010100011111000; end
            14'd15950 : begin out <= 64'b1010100111010101101010101000100100011111100010011010110000000100; end
            14'd15951 : begin out <= 64'b1010101001000010101010001011100000101010101110100010101110100000; end
            14'd15952 : begin out <= 64'b0010011110000000001010011001010110101011101001000001011110000100; end
            14'd15953 : begin out <= 64'b0010000000101101001001011010110100100100111111100010100001001101; end
            14'd15954 : begin out <= 64'b1010011100000010001001011110001100100101001100011010000000000011; end
            14'd15955 : begin out <= 64'b1010010101001100001000110111101010011100001010011010101111101010; end
            14'd15956 : begin out <= 64'b1010010000010100101001010110011100010110111001111010100100110011; end
            14'd15957 : begin out <= 64'b1001111111000100101010110101110010100110010000110010100110011110; end
            14'd15958 : begin out <= 64'b1010100100100101101010001111011110100111100110010010100001101010; end
            14'd15959 : begin out <= 64'b0010100111100101100111101011111000101010001100010010100110100000; end
            14'd15960 : begin out <= 64'b0010100110101000101000001111101110011100101100000010100101100111; end
            14'd15961 : begin out <= 64'b0010101010001111101010000001110100100010101100010010101101010011; end
            14'd15962 : begin out <= 64'b1010001111010000101000100000101100100110011101010010000011010100; end
            14'd15963 : begin out <= 64'b0010101010111011001001111110011000100100111110001010001101111001; end
            14'd15964 : begin out <= 64'b1010000001000001101010101001111000100011101101110010000011100111; end
            14'd15965 : begin out <= 64'b1010101110001100001010001010010110101011111111100010010001101101; end
            14'd15966 : begin out <= 64'b1010100110010001001010010101101100101011011111111010101011001101; end
            14'd15967 : begin out <= 64'b0010100100110001101000010000111100100000001011110010010011011001; end
            14'd15968 : begin out <= 64'b0010000111110110101010101101011000100111001101000010001001100100; end
            14'd15969 : begin out <= 64'b1010101110110110001010001101110110101001001100110001110010010101; end
            14'd15970 : begin out <= 64'b1000111001100000001010111001011010101000010010011010001011010111; end
            14'd15971 : begin out <= 64'b0001111000001100001010000001000110101001011110111001110100000010; end
            14'd15972 : begin out <= 64'b1001011101000001101010010001100100100101011100110010010010111101; end
            14'd15973 : begin out <= 64'b0010010101001011001010000001011000101001011101000010101110011001; end
            14'd15974 : begin out <= 64'b1010101000010001101010001010100110010100010111011010010010000101; end
            14'd15975 : begin out <= 64'b1010010010000010000101011101011100101011011110110010001100011111; end
            14'd15976 : begin out <= 64'b0010001000000000001010110010011000100111110100100010100111000010; end
            14'd15977 : begin out <= 64'b1001110010001111001010010100010110100100010101110010000000000001; end
            14'd15978 : begin out <= 64'b0010001111011100101010010110001000100000100010111010101011001111; end
            14'd15979 : begin out <= 64'b1001100010001110001001010010100000101010111100110001101100110101; end
            14'd15980 : begin out <= 64'b0010100100001001101010111000111010101010011001000001111011111000; end
            14'd15981 : begin out <= 64'b1010100111110101001001101001110110101001100111111010100111001010; end
            14'd15982 : begin out <= 64'b1010100101110001101010100101010010100111101100001010010010011000; end
            14'd15983 : begin out <= 64'b1010011101010100101001101110110110011001010110010010100001110011; end
            14'd15984 : begin out <= 64'b1010100101101011000101111101010010100100010110010010010001011000; end
            14'd15985 : begin out <= 64'b0010101000010111101001001001000110100000110101001010100010001101; end
            14'd15986 : begin out <= 64'b1010011101010101001000001111101010100101101010011010101111010000; end
            14'd15987 : begin out <= 64'b0001110001010110100111010101000110101001000010110010101111000111; end
            14'd15988 : begin out <= 64'b0010100110011100001001011101011000101000011011100010100101000010; end
            14'd15989 : begin out <= 64'b0010100011100000001010001011010110100111010000100010101010100100; end
            14'd15990 : begin out <= 64'b1010101111101011101010000101001010011111001100101010101011011011; end
            14'd15991 : begin out <= 64'b0010000011000000001010011010100010100111101010001010100001110111; end
            14'd15992 : begin out <= 64'b0010101011111011001010110011011100101001011111111010011010011010; end
            14'd15993 : begin out <= 64'b0010101010111000101001111111111010100111110010000010100000010001; end
            14'd15994 : begin out <= 64'b1010000110001111101010101100000010100001100100000010100000011111; end
            14'd15995 : begin out <= 64'b1010100010111101101010111010110000010110100000111010101001101111; end
            14'd15996 : begin out <= 64'b1010010001101011000100110010001000101001111000000010101010010110; end
            14'd15997 : begin out <= 64'b0010001110010011001010001011000110101010000010000001101100011110; end
            14'd15998 : begin out <= 64'b1010000001101110101001001111101010101010111001011010011101010000; end
            14'd15999 : begin out <= 64'b1010100000110100101001110000100000100110010100010010011100011110; end
            14'd16000 : begin out <= 64'b0010001011011101001001111001000010101011010111011010101001111111; end
            14'd16001 : begin out <= 64'b1010011111110000001001011100111000011110000000110010100111001010; end
            14'd16002 : begin out <= 64'b0010100001011110101010111010110000101010111010111000011110001010; end
            14'd16003 : begin out <= 64'b0010000011010101101010010111011010100011111111010010101111011001; end
            14'd16004 : begin out <= 64'b1010010011110101101010110010111010101010011011001010100000001010; end
            14'd16005 : begin out <= 64'b1001110110110111001010110011000010101011011000100010100001100111; end
            14'd16006 : begin out <= 64'b1001111011011010101001111111010100011100101001110010100101111101; end
            14'd16007 : begin out <= 64'b1001100101000011101000100011001000101001110000000010100111010101; end
            14'd16008 : begin out <= 64'b0010011111001011001010000100011110101011010110110010010011010000; end
            14'd16009 : begin out <= 64'b0010011101100000101000010110000010100001010110100010000011001100; end
            14'd16010 : begin out <= 64'b1010011001100110101010010100010000101000001110111010100001011100; end
            14'd16011 : begin out <= 64'b0010100101011010101010101110011000100101100110101010101110101111; end
            14'd16012 : begin out <= 64'b1010010011101110101010001101010100101001011001110010101010001001; end
            14'd16013 : begin out <= 64'b1010100100100110101010001100000000101001011111011000110011110100; end
            14'd16014 : begin out <= 64'b0010101000010000101010000010110000101010100011110010101000000110; end
            14'd16015 : begin out <= 64'b0010100000101010001001010101010000011110000100101010001100101100; end
            14'd16016 : begin out <= 64'b0010011010111100001010000101110000101011111110111001110110111000; end
            14'd16017 : begin out <= 64'b0010101111100010001010010101100110100001010100001000111000111111; end
            14'd16018 : begin out <= 64'b0010100111001010101000011000011000101001000101100010011111001101; end
            14'd16019 : begin out <= 64'b0010100011111110000111011110000000010000010101010010100000011001; end
            14'd16020 : begin out <= 64'b0010101110000101001001110111111000100101111101011010100101101111; end
            14'd16021 : begin out <= 64'b0010001111000110001001011000100000101011001011011001010001010110; end
            14'd16022 : begin out <= 64'b0010101011100010101010101010110010101010101101010010011011101101; end
            14'd16023 : begin out <= 64'b1010010001111011101000011000011100100010100000111010100110110101; end
            14'd16024 : begin out <= 64'b1010011010101001000110001110100000101011010011001001100101110110; end
            14'd16025 : begin out <= 64'b1010011110110111101000011011011100100101110111110010100010101100; end
            14'd16026 : begin out <= 64'b0001111111000011001000111010001110101000100101110010000111100111; end
            14'd16027 : begin out <= 64'b0010010000100101101000110000011110100110101111000010100101011111; end
            14'd16028 : begin out <= 64'b0010100000010011101010011010110100100111001001011010100101110000; end
            14'd16029 : begin out <= 64'b0010100001001100001010010010000010100011101111100010100111000100; end
            14'd16030 : begin out <= 64'b1010010011111000001010101110111110100111010010111001000001111011; end
            14'd16031 : begin out <= 64'b0010101011100101001010011010011000100111110110010010010001111101; end
            14'd16032 : begin out <= 64'b1010010001010101001010101011110010100110010110011001101111010001; end
            14'd16033 : begin out <= 64'b1010101010000000101010011001100110101010001001100010100000000100; end
            14'd16034 : begin out <= 64'b1001111000000111001010000111001100101011111101000010000001000010; end
            14'd16035 : begin out <= 64'b1010100011101010000101000110100010010110011010010010101100000000; end
            14'd16036 : begin out <= 64'b0010100111011000101000011010100110011111110100100010100111011111; end
            14'd16037 : begin out <= 64'b0010010011110110101000100111010110101001111001101001100001000001; end
            14'd16038 : begin out <= 64'b1001110001010110101010110110010000101010111001101000110110110110; end
            14'd16039 : begin out <= 64'b0010010011101110101010001101101100101010101011011010000110000001; end
            14'd16040 : begin out <= 64'b0010100000100111101001101001001010100110101101011010010100101000; end
            14'd16041 : begin out <= 64'b0010010101010110001001101101101000100001000010100010010110110011; end
            14'd16042 : begin out <= 64'b1010010000011000001010110110011110100011101001110010011001101110; end
            14'd16043 : begin out <= 64'b1010011000111001001001011010001100101000001100001010101111000010; end
            14'd16044 : begin out <= 64'b1010100001100100101001100101011000100101001000011010101001101100; end
            14'd16045 : begin out <= 64'b0010000000110100001000001001111110101010010111101010001001000011; end
            14'd16046 : begin out <= 64'b1010010000011110001000110100011010100000100110011010011011101110; end
            14'd16047 : begin out <= 64'b0010011100010000101010101011010100100110010110010010101100101011; end
            14'd16048 : begin out <= 64'b1010000100011010101010111001110100101001101100000010100000000001; end
            14'd16049 : begin out <= 64'b0010011111100101101001010110101100101001101000111010101010111100; end
            14'd16050 : begin out <= 64'b1010011100101011101000011101111000101000000001001010100110010000; end
            14'd16051 : begin out <= 64'b0010000111111100001010101000100010100010110101101001110110110101; end
            14'd16052 : begin out <= 64'b0010100001010011101010110111110010101011111110100010001011011010; end
            14'd16053 : begin out <= 64'b1010101000011010001000001111110110011101011110110010000000110101; end
            14'd16054 : begin out <= 64'b0010001010001011101001001000110110100111101110101010101100001100; end
            14'd16055 : begin out <= 64'b1001110000011110101000100001101010101001011111010001001100011100; end
            14'd16056 : begin out <= 64'b0010011100011001001011000000000010100000011011110010011110011111; end
            14'd16057 : begin out <= 64'b1010010111001001001000011001110010101010001110010010011100101011; end
            14'd16058 : begin out <= 64'b0010100010000110101000000000101110101011111111111010100011111100; end
            14'd16059 : begin out <= 64'b0010100100100001001010100101100000001100110000101010010010000000; end
            14'd16060 : begin out <= 64'b0010100000010111101010010101110010100100011101001010101000001010; end
            14'd16061 : begin out <= 64'b0010100001010000001010110011101010011111011000100010100101011000; end
            14'd16062 : begin out <= 64'b1010101100010101001010001100011110101000110010010010011111101111; end
            14'd16063 : begin out <= 64'b0010101100110011101010001110101010101000001011111010100111111100; end
            14'd16064 : begin out <= 64'b0010000111001101101010011101000100101000001010000010100010101000; end
            14'd16065 : begin out <= 64'b1010101100001100001000110101100110100111000100101010100100101011; end
            14'd16066 : begin out <= 64'b1010100100000011001001011011110100101000000000111010101010001000; end
            14'd16067 : begin out <= 64'b0010001000111010001000010100110000100001111111111010010101111111; end
            14'd16068 : begin out <= 64'b1010000011011111001001011011000010101010010101100010101100010110; end
            14'd16069 : begin out <= 64'b0010101101100001001010001101100100100011010010011001001111111110; end
            14'd16070 : begin out <= 64'b0000100100001011001010110001010010101011111001100010101001000001; end
            14'd16071 : begin out <= 64'b0001101111100110101000000111011010100111010111110010101001000110; end
            14'd16072 : begin out <= 64'b0010100100011111001001010110100110100101101111110010011101000010; end
            14'd16073 : begin out <= 64'b0010011011111011001000011010110010101010010000010010001110100001; end
            14'd16074 : begin out <= 64'b1010101000011011001010111001011100101010000111000010011100001011; end
            14'd16075 : begin out <= 64'b1010100011110010101000100010000110100110010110010010100001000010; end
            14'd16076 : begin out <= 64'b0010010110110110001010100100001010100100110001000010101011011000; end
            14'd16077 : begin out <= 64'b0010010011110111101000100110010110101011000110111001101000101001; end
            14'd16078 : begin out <= 64'b1001010111011100101000111101100000101000100101111010010111111001; end
            14'd16079 : begin out <= 64'b1010101010011110101001110100111000011100001010111010001011000100; end
            14'd16080 : begin out <= 64'b0010101101110001101000110001111000000101000000110010100000010110; end
            14'd16081 : begin out <= 64'b0010101100111111101010000100100100100101111111000010100011111100; end
            14'd16082 : begin out <= 64'b1010011000011000101010111000010000100100001010100010010110100100; end
            14'd16083 : begin out <= 64'b1010001000111000001010100100010110101010101111111010101000001010; end
            14'd16084 : begin out <= 64'b0010001100000101101010100110111110100111011110111010101000111110; end
            14'd16085 : begin out <= 64'b1010101010011101001000011111001110101010101010001010010111100000; end
            14'd16086 : begin out <= 64'b1010101101100001101010010111111100000101011010100010010111111111; end
            14'd16087 : begin out <= 64'b1010000101100111101001010010111100100010111110111010101101001111; end
            14'd16088 : begin out <= 64'b0010010111101100001001000101010100101001011100101010010000100001; end
            14'd16089 : begin out <= 64'b1010100110001110101010100100011000100111010100001010000001110100; end
            14'd16090 : begin out <= 64'b0001101100011011000110111001000010100111010000000001111111111010; end
            14'd16091 : begin out <= 64'b1010100101000010000101000111010100011011111011111010011010111010; end
            14'd16092 : begin out <= 64'b1010100100111000000111111001001010100001111100010010001011000101; end
            14'd16093 : begin out <= 64'b1010011111000111001001000010110000101010110101101010100011101010; end
            14'd16094 : begin out <= 64'b1010100100100011101001111000000110101011110010100010101000010000; end
            14'd16095 : begin out <= 64'b0010100100011111101000001001011010100101001010011010100010101101; end
            14'd16096 : begin out <= 64'b0010100100010010001010101111111110100111110110010010011000100100; end
            14'd16097 : begin out <= 64'b0010100101100110101010010111110100101011110011001010101000111101; end
            14'd16098 : begin out <= 64'b0010100001101100001000011110111100100111010000001001111110110100; end
            14'd16099 : begin out <= 64'b1010101100111000001010011100111000011011001010101010010100001111; end
            14'd16100 : begin out <= 64'b1010101000111100001001011001101010101011011011001010010110010101; end
            14'd16101 : begin out <= 64'b1010011101010001101010001011101100101000011100001010100001010011; end
            14'd16102 : begin out <= 64'b1010100000001000101001011110011000011011101011010010010010010101; end
            14'd16103 : begin out <= 64'b1010101001000000001001100111011110100101100110111010100111110010; end
            14'd16104 : begin out <= 64'b0010001010101000101010000111010110101010011100011010000010110111; end
            14'd16105 : begin out <= 64'b1010001100000100100110001001110110100010000010011010101101100011; end
            14'd16106 : begin out <= 64'b0010001011000101101010101101011000100101010001011001100001000001; end
            14'd16107 : begin out <= 64'b1010101101000001001000111010111000100111110000011010000101000110; end
            14'd16108 : begin out <= 64'b0010101001001100101001010001010110101011011010000001110011000110; end
            14'd16109 : begin out <= 64'b1010100100000100000111011111110000101010101110101010010000010100; end
            14'd16110 : begin out <= 64'b1010000010011001001010000111101000010011110100111001111000010111; end
            14'd16111 : begin out <= 64'b1010101110011000001001101000010000101001100000101010100001111110; end
            14'd16112 : begin out <= 64'b1010100101111000001001001101110100100010010110011001100100110010; end
            14'd16113 : begin out <= 64'b1010100010000101001010100001110100101000011110100010010011101111; end
            14'd16114 : begin out <= 64'b0010100001111000101000100010110010101000001100110010100101011110; end
            14'd16115 : begin out <= 64'b1010010110001000101010001001100000010110001110010010101111010011; end
            14'd16116 : begin out <= 64'b1010100100100000001010111011010100101011011111101010101011101011; end
            14'd16117 : begin out <= 64'b1010000110111000001010011101101010101010101011010010101011111001; end
            14'd16118 : begin out <= 64'b0010011001000000101010000100001100101011110101100010000011011000; end
            14'd16119 : begin out <= 64'b0001001011111100101010000111011010101000100000111010001101101001; end
            14'd16120 : begin out <= 64'b1010101011010100001001000001001100101011000011100010011010000000; end
            14'd16121 : begin out <= 64'b1010001100100011101010111110010010011010010101010010101101000011; end
            14'd16122 : begin out <= 64'b0010100000110100001010101011001010100000111100110001110101101100; end
            14'd16123 : begin out <= 64'b1010010011110101101001000001111100100010100010001010101100001011; end
            14'd16124 : begin out <= 64'b1010100111011000001010011011000100100111001000000010101100001000; end
            14'd16125 : begin out <= 64'b1010100000000101101010000111000000100111000011100010100001011101; end
            14'd16126 : begin out <= 64'b0010011110101100101001110100110100100111000011101010101101100110; end
            14'd16127 : begin out <= 64'b0001100100100100001010000011011110101011101000111010100011111111; end
            14'd16128 : begin out <= 64'b1010010001111010001010111111010110100110110000011010011011001101; end
            14'd16129 : begin out <= 64'b0010100110000010101010100000000000100100001100110010100111000011; end
            14'd16130 : begin out <= 64'b1010101110011111101001000011011100100111001111011010100000110111; end
            14'd16131 : begin out <= 64'b1010101000100001101000001101011100011011011011101010010000110101; end
            14'd16132 : begin out <= 64'b0010100001010010001010001111001000100011101111110010010111111011; end
            14'd16133 : begin out <= 64'b0010011101010000001010011110110110011111000101110010010011001011; end
            14'd16134 : begin out <= 64'b1010100100111111001010001100000000101000001101111010001011100101; end
            14'd16135 : begin out <= 64'b1010100111101010001010101000011110100101010101100010000110000001; end
            14'd16136 : begin out <= 64'b1010101000100100001010010101101100101001110011001010100110100100; end
            14'd16137 : begin out <= 64'b0010101111000101101010101101000100101001000000111010000001100100; end
            14'd16138 : begin out <= 64'b0010100011110110101000001100101100011110110100011010100111001101; end
            14'd16139 : begin out <= 64'b0010100110011010001010110101001010100101110101000010101011101010; end
            14'd16140 : begin out <= 64'b1010101000001101001001101100011110101000010001100010100001101001; end
            14'd16141 : begin out <= 64'b1010001110101000001000100111000000011000101100111001011100010011; end
            14'd16142 : begin out <= 64'b1010010110000110101001101001010100101011001011111000101111111011; end
            14'd16143 : begin out <= 64'b1010101001101000101010001011010010100000010101010010001110101011; end
            14'd16144 : begin out <= 64'b1010010001111000001000110110010000100111110100110010100010011111; end
            14'd16145 : begin out <= 64'b1010100111010000001001001110110100100010010001100010011011010100; end
            14'd16146 : begin out <= 64'b0010010110101011001010101100111100100010010011001010101111001000; end
            14'd16147 : begin out <= 64'b0010010100001110101010100010110100101000010100011010011101100110; end
            14'd16148 : begin out <= 64'b1010100101010001001010110001110010101000000111010010101000101101; end
            14'd16149 : begin out <= 64'b1010101010101110001010101000110110100101111011100010010100011011; end
            14'd16150 : begin out <= 64'b0010101000010101001010100100011110100101001100110010100111001010; end
            14'd16151 : begin out <= 64'b0010101110000100001001011100000110100100000001110010010000110111; end
            14'd16152 : begin out <= 64'b0010010011111101100111001001010010100100001000100010011101110010; end
            14'd16153 : begin out <= 64'b0010011111100000000111101110001010101010110001011010010101111110; end
            14'd16154 : begin out <= 64'b1010001110100111001011000001001100100111100101111010100100011001; end
            14'd16155 : begin out <= 64'b1010011010100101101001000000010000100111111011111010101100000100; end
            14'd16156 : begin out <= 64'b1010101010010101100100110000001010011000100111000010010010001100; end
            14'd16157 : begin out <= 64'b0010001110100001001000000001001000101001100100001010101111010110; end
            14'd16158 : begin out <= 64'b0010010100110010101001101111000110101011010101000010101110001011; end
            14'd16159 : begin out <= 64'b1010001110101100101010110110001010101011001100010010010100000101; end
            14'd16160 : begin out <= 64'b0001011001111110001010000110101110101010111111000010100100010111; end
            14'd16161 : begin out <= 64'b0010100001010101101010010111010100100101100001100010101110101000; end
            14'd16162 : begin out <= 64'b0010101011100111101010111100101100101000111101011010100101110111; end
            14'd16163 : begin out <= 64'b0010010111011001101001010000001010100110001101101010100100110010; end
            14'd16164 : begin out <= 64'b0010011011110101001010100111001100101010011111101010100111101110; end
            14'd16165 : begin out <= 64'b1010101001111000001010000001011100101001100110010010100111100100; end
            14'd16166 : begin out <= 64'b1001100010011100001010101001011000101010100010101010101101100111; end
            14'd16167 : begin out <= 64'b0001111100011100001010111111111000101011010111011001011011100101; end
            14'd16168 : begin out <= 64'b0010100010100011101010110101111000100011000111110010101111110000; end
            14'd16169 : begin out <= 64'b1010010011110000101010001001010010101010001101100010100100100010; end
            14'd16170 : begin out <= 64'b1001101101011111001001011100111000101001011000111001111111100110; end
            14'd16171 : begin out <= 64'b1010100100101000101001110101000110101010011010011010101101110110; end
            14'd16172 : begin out <= 64'b1010100111010111001010000010000010101001110111001010100010110010; end
            14'd16173 : begin out <= 64'b1010101011111110101010001110100110100100011001000010010011100101; end
            14'd16174 : begin out <= 64'b1010010100100110101001110111110010011110001101101010011110101000; end
            14'd16175 : begin out <= 64'b1010010110101101001001011000101010101011100110000010101000100110; end
            14'd16176 : begin out <= 64'b1010100111101110001010101000111000100101101001111010010001011110; end
            14'd16177 : begin out <= 64'b1010100100110100001001100000001000100110110000001010101111001011; end
            14'd16178 : begin out <= 64'b0010101100010001001001101110100010100101010111000010100011000000; end
            14'd16179 : begin out <= 64'b1010010010011010001001001000101100011100101001010010101000000110; end
            14'd16180 : begin out <= 64'b1010101000110110000110010101000000100100000000000010101101100111; end
            14'd16181 : begin out <= 64'b0010101100001111001010111100011000100011110101111010010001101001; end
            14'd16182 : begin out <= 64'b1010011100000100101010001101110000100111011101000010101101101101; end
            14'd16183 : begin out <= 64'b0010101011101110101010111110010100101000011110100010100001001001; end
            14'd16184 : begin out <= 64'b1010100001110101101010111101001110101000100011001010011011011111; end
            14'd16185 : begin out <= 64'b1010001110100101101010100100010110101010011100101010101010010011; end
            14'd16186 : begin out <= 64'b1010100100100111101001011101001000100101101111101010010011101110; end
            14'd16187 : begin out <= 64'b1010101111010010001001001110001010100110010100111010100011100111; end
            14'd16188 : begin out <= 64'b0010100001100100000111001011101000010111001100010010000011011100; end
            14'd16189 : begin out <= 64'b1001110110011001001010010011110100101001100110100010011000100101; end
            14'd16190 : begin out <= 64'b0010010110110010001000110011001100101011101010011010000100000111; end
            14'd16191 : begin out <= 64'b1010100010110001101010000101111110101010110111110001111111000001; end
            14'd16192 : begin out <= 64'b1010010011010011001001011101100100100000001001101010011010101010; end
            14'd16193 : begin out <= 64'b0010011000111000100111001010001110101011000111001010010001011110; end
            14'd16194 : begin out <= 64'b0001101011001100001010111010010010100101110010111010010111001011; end
            14'd16195 : begin out <= 64'b0010010101101000000111110110100110100100010101110010101101111111; end
            14'd16196 : begin out <= 64'b1010100111010110101010001010100100100000010011100010101110011101; end
            14'd16197 : begin out <= 64'b1001010101000101101010110010110100100011001010111010011101000011; end
            14'd16198 : begin out <= 64'b1010000010100110101000110111101110100001011100010010010101110111; end
            14'd16199 : begin out <= 64'b1010100101011101001001101001101110100111100011011001111111010101; end
            14'd16200 : begin out <= 64'b0010101100100100001001011100010000101011011111100010001010101111; end
            14'd16201 : begin out <= 64'b0010100101101001101011000001001110101010010011100010101010010010; end
            14'd16202 : begin out <= 64'b1010100000101111001001000000001010100010110100100010101010011101; end
            14'd16203 : begin out <= 64'b1010011111101111001001000001000010100000001000110010011110000001; end
            14'd16204 : begin out <= 64'b1010001001000101101010001100000100100000101010010010101100010001; end
            14'd16205 : begin out <= 64'b1010101101000001001000000101010000101000001110001010101010010110; end
            14'd16206 : begin out <= 64'b1010100101000001001010100110010000100111011011000001111011011101; end
            14'd16207 : begin out <= 64'b1010010100100111101001101000011000100110000010011010000101001010; end
            14'd16208 : begin out <= 64'b0000000100001010101010010001110010101001010100100010101111000001; end
            14'd16209 : begin out <= 64'b0010100000011000000111011000000100100100000101110010010000100011; end
            14'd16210 : begin out <= 64'b1010101010100100101010010010111110101001110011010000110110110110; end
            14'd16211 : begin out <= 64'b1010000110010001101010100011110000101010001110111010101100111011; end
            14'd16212 : begin out <= 64'b1010011100111010001010111100001100100001101111010001101001010100; end
            14'd16213 : begin out <= 64'b0010100101111101000101011000000110100001101011010010000101101011; end
            14'd16214 : begin out <= 64'b0010101000000101101010011010100100101010001000010010100100011001; end
            14'd16215 : begin out <= 64'b1010001001110011101010111011101000101010001010011001110100001100; end
            14'd16216 : begin out <= 64'b1010100010100100101010000100010110101001010111011010100011010001; end
            14'd16217 : begin out <= 64'b0001100100111010101001110001010100101001111010011010101011101000; end
            14'd16218 : begin out <= 64'b0010101000001011101010000100010010101000001101010010011010000101; end
            14'd16219 : begin out <= 64'b0010011111000100101001000111111000101011100101010010101010010110; end
            14'd16220 : begin out <= 64'b1010010001011100101010000010110100101010000000010010100001011111; end
            14'd16221 : begin out <= 64'b0010101000000010101010111101111000101011111110111010100100010000; end
            14'd16222 : begin out <= 64'b0010100100001101001010111011100110011110011001010010100011001110; end
            14'd16223 : begin out <= 64'b0010101001110101101010101000111010100000000110010010100101110111; end
            14'd16224 : begin out <= 64'b1010010100110001001000001000001100011110001111111000111010110100; end
            14'd16225 : begin out <= 64'b0010011011101001100111001101111000100011110101111001111001011011; end
            14'd16226 : begin out <= 64'b0010100010110100101001011110000010100001100100010010101000000001; end
            14'd16227 : begin out <= 64'b1010101000111010101010000110111010101011110001011010010010110101; end
            14'd16228 : begin out <= 64'b1010101001100011000101100111000000011000111010001010000010100000; end
            14'd16229 : begin out <= 64'b1010000000111010001010110010110010101000000101110010101010100100; end
            14'd16230 : begin out <= 64'b0010010010100000100101101011111110101010001000101010101011111010; end
            14'd16231 : begin out <= 64'b1010101111001101000111001100111010101010000001111001111010000111; end
            14'd16232 : begin out <= 64'b1010010000011101001010001111001000101010000011110010101001011000; end
            14'd16233 : begin out <= 64'b1010101110101010001001111101011000101000011111011010010010101111; end
            14'd16234 : begin out <= 64'b0010101111000001001001011101100010101010110110110010000000111000; end
            14'd16235 : begin out <= 64'b1010101000011010101010101101011000101011101101011010000110011010; end
            14'd16236 : begin out <= 64'b0010101010000110001001011011110000011110101100111001101011101000; end
            14'd16237 : begin out <= 64'b0010011000100101001010001101111000101001010010100010100001000111; end
            14'd16238 : begin out <= 64'b1010011110101111001010111000000110100001011011110010100111011111; end
            14'd16239 : begin out <= 64'b1010011011111011101010000110011110100000010101101010011010000111; end
            14'd16240 : begin out <= 64'b0010010000001101001000010111010000011000110110110001101000001001; end
            14'd16241 : begin out <= 64'b0010011010010111100100011000010100100101000000010010101101001011; end
            14'd16242 : begin out <= 64'b0010101110000111100110100010110100011111001011001010001100101000; end
            14'd16243 : begin out <= 64'b1010010100100100001010100001110000101010011100100010010000001000; end
            14'd16244 : begin out <= 64'b0010100100110101001010101111000000100101110100000010011100100010; end
            14'd16245 : begin out <= 64'b1001110001100000101001101000101000100101100010000010101101111111; end
            14'd16246 : begin out <= 64'b1001111000100111101010000110111010100100111111010010101101111101; end
            14'd16247 : begin out <= 64'b0001101101111001001000101001100010100100100111110010010010100000; end
            14'd16248 : begin out <= 64'b1001111111100010001001011100101010101011001110101010100000111010; end
            14'd16249 : begin out <= 64'b0010010100101100001000101000110010101000111111101010000001000001; end
            14'd16250 : begin out <= 64'b0001101010111110001010110001101110101011110110111010011001110110; end
            14'd16251 : begin out <= 64'b1010100101010110101000111011011100101100000000000010101101011000; end
            14'd16252 : begin out <= 64'b0010101001111110101010011000101100100101110100001010010101110100; end
            14'd16253 : begin out <= 64'b1010100111001001101001011110101100101010001001001010101001000001; end
            14'd16254 : begin out <= 64'b1010000100001000000011111101000100101010001110000000100010100011; end
            14'd16255 : begin out <= 64'b0010110000001010001000000110001010101010001011000010101000111110; end
            14'd16256 : begin out <= 64'b0010001101101101001010000010000010011100111110001010101100010011; end
            14'd16257 : begin out <= 64'b1001111010110101101001101010110000101011000100010001011000100011; end
            14'd16258 : begin out <= 64'b0010101111100100101010101011001100100110110111111010100000110011; end
            14'd16259 : begin out <= 64'b1010010100111010101010000001000010101001011101111010101110101100; end
            14'd16260 : begin out <= 64'b0010010011001100001010000011101000100111111110001010010000000101; end
            14'd16261 : begin out <= 64'b1010100111010101101001110110000110100011001001000010101000010110; end
            14'd16262 : begin out <= 64'b0010101010110110101001111011010010101010111100100010100100001001; end
            14'd16263 : begin out <= 64'b0010100101100101001001001100011000101011011001010001110110111000; end
            14'd16264 : begin out <= 64'b1010011100010100101001110001110100100110011011000010100001100010; end
            14'd16265 : begin out <= 64'b1001011110010011001010100010000000101010001111110010100000110100; end
            14'd16266 : begin out <= 64'b1010010001111010001010001011011010100101101000000010100010011001; end
            14'd16267 : begin out <= 64'b0010011111001001101000110111010000100111001110011010100001001110; end
            14'd16268 : begin out <= 64'b0010101001000011101001101010100110101000010001011010000010000011; end
            14'd16269 : begin out <= 64'b1010001101110100001010000111000010101011011101000010001111010000; end
            14'd16270 : begin out <= 64'b1001111110001111101010011110101010101010110100000010011101110000; end
            14'd16271 : begin out <= 64'b0010100110110010101010010000011000101000100100101010010000010001; end
            14'd16272 : begin out <= 64'b0010001000010110101000111110101100100100010010111001111101000001; end
            14'd16273 : begin out <= 64'b1010100110011000001010000000000010011101100010010010010100011010; end
            14'd16274 : begin out <= 64'b0010100000111110101010001000011100101001101010000010100100000111; end
            14'd16275 : begin out <= 64'b1010010100100101101001111110101000101010101000111010100100111010; end
            14'd16276 : begin out <= 64'b0001101010011110001001101001010100101000001101111010100000101111; end
            14'd16277 : begin out <= 64'b0010010001110111001000111010101000011000110000010010101000001110; end
            14'd16278 : begin out <= 64'b0010100111100001101000010011011100100110011101101010011100011000; end
            14'd16279 : begin out <= 64'b0010100111110101001010001010110100101000001011111010101111101101; end
            14'd16280 : begin out <= 64'b1001110000010110000011101011011010101011001100000010100000010000; end
            14'd16281 : begin out <= 64'b1010010101011100001010000101100010011100100000101010011111111001; end
            14'd16282 : begin out <= 64'b1010100101110011000110010001001110011100001000011010010110111010; end
            14'd16283 : begin out <= 64'b1010100111100010101001110010101110101010110110010010101100110011; end
            14'd16284 : begin out <= 64'b0010011000101100101010101010110000101001000011000010011101111101; end
            14'd16285 : begin out <= 64'b1000111110000100101010000010111000100110000011010010101111011010; end
            14'd16286 : begin out <= 64'b1010110000001010101010011011101110100110100011111001111001011100; end
            14'd16287 : begin out <= 64'b1001101010111111001001101000111000100110010001101010001101110010; end
            14'd16288 : begin out <= 64'b0001110001010000101001010100001000100100000000111010001100010000; end
            14'd16289 : begin out <= 64'b1001101000011100101010000011011110101001111000001010100000011100; end
            14'd16290 : begin out <= 64'b1010001010001001101000000111000100100000100010110010101001111100; end
            14'd16291 : begin out <= 64'b1010101000001000101010011000110010011100011000011010100101110000; end
            14'd16292 : begin out <= 64'b0010101100111010100111010100111110100100001000100010101110100100; end
            14'd16293 : begin out <= 64'b1010100010111010101010100101000010100001010000101010101110101110; end
            14'd16294 : begin out <= 64'b0010000101111001001000100000001000100101101111011010100111010101; end
            14'd16295 : begin out <= 64'b1010100111011010101001011001001100101001010001010010100010001110; end
            14'd16296 : begin out <= 64'b0001000110001011000111100101100100100011101100110010010111100011; end
            14'd16297 : begin out <= 64'b1010101011100111101000010011101010100011010100000001111100010110; end
            14'd16298 : begin out <= 64'b1010100011000010001010110110111010101001010011000010100000101010; end
            14'd16299 : begin out <= 64'b0010011000010000001010011010101010100110010110101010010111010111; end
            14'd16300 : begin out <= 64'b0010011110010000101010010101111100100100000111110010100000011101; end
            14'd16301 : begin out <= 64'b0010010101011010101010110001011110100110011001001010101010000110; end
            14'd16302 : begin out <= 64'b0001100110011100100111010101011100100111001010101010101001111111; end
            14'd16303 : begin out <= 64'b1010101100001111101010001111010110011100011101011010100110010001; end
            14'd16304 : begin out <= 64'b0010100011010110001010010110111000101001001000101010100010011100; end
            14'd16305 : begin out <= 64'b0010100111100011001000001011010100100101100000111010100000100010; end
            14'd16306 : begin out <= 64'b1001110101110011001010111110111000101010101001011010100011001001; end
            14'd16307 : begin out <= 64'b0010101111001101101001110111110100011010000100101010010111011010; end
            14'd16308 : begin out <= 64'b0010011001001001001010011111110110100110010101011010100111101101; end
            14'd16309 : begin out <= 64'b1010100100000000001010001110110000101000110110001010101111010011; end
            14'd16310 : begin out <= 64'b1001110000011100001010111100111110101010110010001010010011111001; end
            14'd16311 : begin out <= 64'b1010101101000101000110010011010100101000110101010010101000001010; end
            14'd16312 : begin out <= 64'b0010101110001011101010110111010100101000110000001010100011010010; end
            14'd16313 : begin out <= 64'b0010100010011111000111010110000100001101101001101010100010000101; end
            14'd16314 : begin out <= 64'b1001110100100010001010101101100000100100010011000010010001101001; end
            14'd16315 : begin out <= 64'b1010101100110111001010101111010000011001100101111010100111111001; end
            14'd16316 : begin out <= 64'b0010011100000101101010100011010010100011011111101010100000111111; end
            14'd16317 : begin out <= 64'b1010000001111111001010010000001000100111001101101010001010011111; end
            14'd16318 : begin out <= 64'b0010011010101000101001111110011010100011000100101010101011100100; end
            14'd16319 : begin out <= 64'b0001011111000110000011011100110110101011011100100010101000001101; end
            14'd16320 : begin out <= 64'b0010010101011110101010000000010010101011101010101010101110111011; end
            14'd16321 : begin out <= 64'b0010010000011001001010001010100010100110011000111010000011110111; end
            14'd16322 : begin out <= 64'b1010001011100011001001010101100010101001010011111010100111010001; end
            14'd16323 : begin out <= 64'b0000010010110111001010010101100100011000101101000010101100101100; end
            14'd16324 : begin out <= 64'b1010100111110100001010001101011100100100000011110010101101001001; end
            14'd16325 : begin out <= 64'b0010011110100111001010100111101100100110011001100010000010011011; end
            14'd16326 : begin out <= 64'b1010101010110101001010000100010110101011010111010010010011100101; end
            14'd16327 : begin out <= 64'b1010100011000111101010101100011100011000101000100010001110001000; end
            14'd16328 : begin out <= 64'b1010100110000110101010100010011110100100101011000010101011011001; end
            14'd16329 : begin out <= 64'b0010100110101010001010000110100010101010000001101010101110100101; end
            14'd16330 : begin out <= 64'b0010100011010100101010010010101110101011100100011010010000000101; end
            14'd16331 : begin out <= 64'b0010000110000000000111010011110010101000011101100010011000110110; end
            14'd16332 : begin out <= 64'b1010010001001111101000101100100010101000010010100010011011101111; end
            14'd16333 : begin out <= 64'b1010101011000001100110011011110010100111111011111010101011110101; end
            14'd16334 : begin out <= 64'b0010001111000001001010011100111110100111011000100010100110111100; end
            14'd16335 : begin out <= 64'b1001101100100001101010010000110010101001011100001010101000111011; end
            14'd16336 : begin out <= 64'b0010101000001111001001111001000100101001010010101010000111000011; end
            14'd16337 : begin out <= 64'b1010101101011010001001100001110110101001101001101010100001110100; end
            14'd16338 : begin out <= 64'b1010101010010101101010110111111110100010011010111010010100001001; end
            14'd16339 : begin out <= 64'b1001011111101001101000011000001000101000010010011001110010100110; end
            14'd16340 : begin out <= 64'b1010010011101001001010101011100100101001111101001010100100000111; end
            14'd16341 : begin out <= 64'b0010100110000100101010101110110100101000100011010010011000001001; end
            14'd16342 : begin out <= 64'b1010011000011101001010001111111000100010111001000010101110001001; end
            14'd16343 : begin out <= 64'b0010101111001101001000110110100010100011010001111010101000011010; end
            14'd16344 : begin out <= 64'b0010101011110101001000100000010010100101111010001010001010011100; end
            14'd16345 : begin out <= 64'b1010101010100110001010000001100010101011010001101010101011000010; end
            14'd16346 : begin out <= 64'b1010010101111001101000100110100000101000001110011010011101000010; end
            14'd16347 : begin out <= 64'b1010100011101101101000110000111100101000011010111010011010010011; end
            14'd16348 : begin out <= 64'b1001100100111010101010000100100010100111110110100010000101001000; end
            14'd16349 : begin out <= 64'b0010100000111010101010000111010100100101001110110010000111111110; end
            14'd16350 : begin out <= 64'b0001110101010011101000010101110010011111101101010010101010011101; end
            14'd16351 : begin out <= 64'b0010011011111111101010100101101100100100001001000010100100000011; end
            14'd16352 : begin out <= 64'b0010100010101100001000000001000000101001011000010001101010111000; end
            14'd16353 : begin out <= 64'b1010101000011001001010011101000010011111101011011010010010101110; end
            14'd16354 : begin out <= 64'b1010101011101001001001010100000010011110111101110010001000100110; end
            14'd16355 : begin out <= 64'b1010101101000101101010001000011100101000011101110010010010101111; end
            14'd16356 : begin out <= 64'b0010110000010000001001111000100010100100110101000001010000110011; end
            14'd16357 : begin out <= 64'b0010010100001101001001011010011110100101101101110001111000101111; end
            14'd16358 : begin out <= 64'b1010011101111000101001010101110100100101101011111010101100000110; end
            14'd16359 : begin out <= 64'b0001110011110111100101111110101100101000111010010010011011110010; end
            14'd16360 : begin out <= 64'b0010000111010110100110101010110000100111101010011010100101111111; end
            14'd16361 : begin out <= 64'b1001101101110111101001011011101100011101100010111010001100101010; end
            14'd16362 : begin out <= 64'b1010010000110101101011000001010010100001011110101010101011000001; end
            14'd16363 : begin out <= 64'b0010010001001110001010010111001100101001101101001010101111100010; end
            14'd16364 : begin out <= 64'b0001110000010101001010001101001000101000110111111010011110000111; end
            14'd16365 : begin out <= 64'b0010000001011101101000001010001110101010011110111010010110111110; end
            14'd16366 : begin out <= 64'b1010100000000000001010001100101100101010101110100010010010110001; end
            14'd16367 : begin out <= 64'b0000110010100001001000001111011000101001111100111010101011110001; end
            14'd16368 : begin out <= 64'b1010100010101100001010110010010010011010111011000010100011001000; end
            14'd16369 : begin out <= 64'b1010000110101000001010010100110010101010010101010010011101001100; end
            14'd16370 : begin out <= 64'b0010001111010111101010100011101110101000000111001010101100001001; end
            14'd16371 : begin out <= 64'b1010101111100101001001000001001010101000101011000010101010001010; end
            14'd16372 : begin out <= 64'b1010101100000110101010100100001000011001110101100010101111000101; end
            14'd16373 : begin out <= 64'b1001110011110111101001000010101000101010111100000010100111101101; end
            14'd16374 : begin out <= 64'b0010101011001110101001000011010000101011011110001010011010010110; end
            14'd16375 : begin out <= 64'b1010100011001101001000000111000000101000010000111010100001001100; end
            14'd16376 : begin out <= 64'b0010101010001110000111010110011000011110110100100010101101111001; end
            14'd16377 : begin out <= 64'b1010000111100101001001101000010000101001001001000001001101011001; end
            14'd16378 : begin out <= 64'b0010101101111001001001101100011100101010111011101010100110101010; end
            14'd16379 : begin out <= 64'b1010100001000110101010111100111010101001100100110010010100011101; end
            14'd16380 : begin out <= 64'b0010010000101100001010000101110010101000011111110010010011010000; end
            14'd16381 : begin out <= 64'b1010011101011010001010010011001110101010000011110010100101000101; end
            14'd16382 : begin out <= 64'b1010100101110100101000011110000010101000000010001010101110011011; end
            14'd16383 : begin out <= 64'b0010001001101101101010011101111110000010010101010010011011111100; end

        endcase
    end
end
assign data = out;

endmodule //gemm2B
